`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.01.2026 10:08:04
// Design Name: 
// Module Name: Main2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Main2(
    input clk,rst,
    output reg [31:0]sum
    );
    parameter size=137;
    
    reg [size-1:0]ram[size-1:0];
    reg [size-1:0]sumram[size-1:0];
    initial
    begin
        ram[0][0]=1;ram[0][1]=1;ram[0][2]=0;ram[0][3]=1;ram[0][4]=1;ram[0][5]=1;ram[0][6]=1;ram[0][7]=0;ram[0][8]=0;ram[0][9]=1;ram[0][10]=1;ram[0][11]=1;ram[0][12]=0;ram[0][13]=0;ram[0][14]=1;ram[0][15]=1;ram[0][16]=1;ram[0][17]=0;ram[0][18]=1;ram[0][19]=1;ram[0][20]=0;ram[0][21]=1;ram[0][22]=1;ram[0][23]=1;ram[0][24]=1;ram[0][25]=1;ram[0][26]=1;ram[0][27]=1;ram[0][28]=0;ram[0][29]=1;ram[0][30]=1;ram[0][31]=1;ram[0][32]=0;ram[0][33]=1;ram[0][34]=1;ram[0][35]=1;ram[0][36]=1;ram[0][37]=1;ram[0][38]=1;ram[0][39]=1;ram[0][40]=1;ram[0][41]=0;ram[0][42]=1;ram[0][43]=1;ram[0][44]=1;ram[0][45]=1;ram[0][46]=1;ram[0][47]=1;ram[0][48]=1;ram[0][49]=0;ram[0][50]=0;ram[0][51]=1;ram[0][52]=1;ram[0][53]=1;ram[0][54]=1;ram[0][55]=1;ram[0][56]=1;ram[0][57]=0;ram[0][58]=1;ram[0][59]=1;ram[0][60]=0;ram[0][61]=0;ram[0][62]=0;ram[0][63]=0;ram[0][64]=0;ram[0][65]=1;ram[0][66]=1;ram[0][67]=0;ram[0][68]=1;ram[0][69]=0;ram[0][70]=0;ram[0][71]=1;ram[0][72]=0;ram[0][73]=1;ram[0][74]=1;ram[0][75]=1;ram[0][76]=0;ram[0][77]=1;ram[0][78]=0;ram[0][79]=1;ram[0][80]=0;ram[0][81]=1;ram[0][82]=1;ram[0][83]=1;ram[0][84]=0;ram[0][85]=1;ram[0][86]=0;ram[0][87]=0;ram[0][88]=0;ram[0][89]=1;ram[0][90]=1;ram[0][91]=1;ram[0][92]=1;ram[0][93]=1;ram[0][94]=0;ram[0][95]=1;ram[0][96]=0;ram[0][97]=1;ram[0][98]=0;ram[0][99]=1;ram[0][100]=0;ram[0][101]=1;ram[0][102]=0;ram[0][103]=1;ram[0][104]=1;ram[0][105]=1;ram[0][106]=1;ram[0][107]=1;ram[0][108]=1;ram[0][109]=1;ram[0][110]=0;ram[0][111]=0;ram[0][112]=0;ram[0][113]=1;ram[0][114]=0;ram[0][115]=0;ram[0][116]=0;ram[0][117]=1;ram[0][118]=0;ram[0][119]=1;ram[0][120]=0;ram[0][121]=0;ram[0][122]=0;ram[0][123]=1;ram[0][124]=0;ram[0][125]=1;ram[0][126]=0;ram[0][127]=1;ram[0][128]=1;ram[0][129]=1;ram[0][130]=1;ram[0][131]=1;ram[0][132]=1;ram[0][133]=1;ram[0][134]=1;ram[0][135]=1;ram[0][136]=1;
        ram[1][0]=0;ram[1][1]=1;ram[1][2]=0;ram[1][3]=1;ram[1][4]=1;ram[1][5]=0;ram[1][6]=1;ram[1][7]=1;ram[1][8]=0;ram[1][9]=0;ram[1][10]=1;ram[1][11]=1;ram[1][12]=1;ram[1][13]=1;ram[1][14]=1;ram[1][15]=0;ram[1][16]=1;ram[1][17]=0;ram[1][18]=0;ram[1][19]=1;ram[1][20]=0;ram[1][21]=0;ram[1][22]=1;ram[1][23]=1;ram[1][24]=0;ram[1][25]=0;ram[1][26]=1;ram[1][27]=1;ram[1][28]=0;ram[1][29]=1;ram[1][30]=1;ram[1][31]=1;ram[1][32]=0;ram[1][33]=1;ram[1][34]=1;ram[1][35]=0;ram[1][36]=0;ram[1][37]=0;ram[1][38]=1;ram[1][39]=1;ram[1][40]=0;ram[1][41]=1;ram[1][42]=0;ram[1][43]=1;ram[1][44]=0;ram[1][45]=1;ram[1][46]=0;ram[1][47]=1;ram[1][48]=0;ram[1][49]=0;ram[1][50]=1;ram[1][51]=0;ram[1][52]=0;ram[1][53]=1;ram[1][54]=1;ram[1][55]=0;ram[1][56]=1;ram[1][57]=1;ram[1][58]=1;ram[1][59]=1;ram[1][60]=0;ram[1][61]=1;ram[1][62]=0;ram[1][63]=1;ram[1][64]=1;ram[1][65]=1;ram[1][66]=1;ram[1][67]=1;ram[1][68]=1;ram[1][69]=1;ram[1][70]=1;ram[1][71]=0;ram[1][72]=1;ram[1][73]=1;ram[1][74]=0;ram[1][75]=1;ram[1][76]=0;ram[1][77]=1;ram[1][78]=0;ram[1][79]=1;ram[1][80]=0;ram[1][81]=1;ram[1][82]=1;ram[1][83]=1;ram[1][84]=0;ram[1][85]=0;ram[1][86]=1;ram[1][87]=1;ram[1][88]=1;ram[1][89]=1;ram[1][90]=1;ram[1][91]=0;ram[1][92]=0;ram[1][93]=1;ram[1][94]=0;ram[1][95]=1;ram[1][96]=1;ram[1][97]=1;ram[1][98]=0;ram[1][99]=1;ram[1][100]=0;ram[1][101]=1;ram[1][102]=0;ram[1][103]=0;ram[1][104]=1;ram[1][105]=1;ram[1][106]=0;ram[1][107]=0;ram[1][108]=1;ram[1][109]=1;ram[1][110]=0;ram[1][111]=1;ram[1][112]=1;ram[1][113]=1;ram[1][114]=0;ram[1][115]=1;ram[1][116]=0;ram[1][117]=0;ram[1][118]=0;ram[1][119]=1;ram[1][120]=1;ram[1][121]=0;ram[1][122]=1;ram[1][123]=1;ram[1][124]=1;ram[1][125]=1;ram[1][126]=1;ram[1][127]=0;ram[1][128]=1;ram[1][129]=0;ram[1][130]=0;ram[1][131]=1;ram[1][132]=0;ram[1][133]=0;ram[1][134]=1;ram[1][135]=0;ram[1][136]=1;
        ram[2][0]=0;ram[2][1]=1;ram[2][2]=0;ram[2][3]=1;ram[2][4]=1;ram[2][5]=1;ram[2][6]=0;ram[2][7]=1;ram[2][8]=1;ram[2][9]=0;ram[2][10]=1;ram[2][11]=0;ram[2][12]=1;ram[2][13]=1;ram[2][14]=0;ram[2][15]=1;ram[2][16]=1;ram[2][17]=1;ram[2][18]=1;ram[2][19]=1;ram[2][20]=0;ram[2][21]=1;ram[2][22]=0;ram[2][23]=1;ram[2][24]=1;ram[2][25]=1;ram[2][26]=0;ram[2][27]=1;ram[2][28]=0;ram[2][29]=1;ram[2][30]=1;ram[2][31]=1;ram[2][32]=1;ram[2][33]=1;ram[2][34]=0;ram[2][35]=1;ram[2][36]=0;ram[2][37]=0;ram[2][38]=0;ram[2][39]=1;ram[2][40]=1;ram[2][41]=1;ram[2][42]=1;ram[2][43]=1;ram[2][44]=1;ram[2][45]=1;ram[2][46]=1;ram[2][47]=1;ram[2][48]=0;ram[2][49]=1;ram[2][50]=1;ram[2][51]=1;ram[2][52]=0;ram[2][53]=1;ram[2][54]=1;ram[2][55]=0;ram[2][56]=1;ram[2][57]=1;ram[2][58]=0;ram[2][59]=1;ram[2][60]=0;ram[2][61]=0;ram[2][62]=1;ram[2][63]=1;ram[2][64]=0;ram[2][65]=0;ram[2][66]=1;ram[2][67]=0;ram[2][68]=1;ram[2][69]=1;ram[2][70]=1;ram[2][71]=1;ram[2][72]=0;ram[2][73]=0;ram[2][74]=1;ram[2][75]=1;ram[2][76]=1;ram[2][77]=0;ram[2][78]=0;ram[2][79]=0;ram[2][80]=1;ram[2][81]=0;ram[2][82]=1;ram[2][83]=0;ram[2][84]=1;ram[2][85]=1;ram[2][86]=1;ram[2][87]=1;ram[2][88]=0;ram[2][89]=0;ram[2][90]=1;ram[2][91]=0;ram[2][92]=0;ram[2][93]=1;ram[2][94]=1;ram[2][95]=0;ram[2][96]=1;ram[2][97]=1;ram[2][98]=0;ram[2][99]=0;ram[2][100]=0;ram[2][101]=1;ram[2][102]=0;ram[2][103]=1;ram[2][104]=0;ram[2][105]=0;ram[2][106]=1;ram[2][107]=1;ram[2][108]=1;ram[2][109]=1;ram[2][110]=1;ram[2][111]=1;ram[2][112]=1;ram[2][113]=0;ram[2][114]=1;ram[2][115]=1;ram[2][116]=1;ram[2][117]=0;ram[2][118]=0;ram[2][119]=1;ram[2][120]=1;ram[2][121]=1;ram[2][122]=0;ram[2][123]=0;ram[2][124]=1;ram[2][125]=1;ram[2][126]=1;ram[2][127]=1;ram[2][128]=0;ram[2][129]=1;ram[2][130]=1;ram[2][131]=1;ram[2][132]=0;ram[2][133]=1;ram[2][134]=1;ram[2][135]=1;ram[2][136]=1;
        ram[3][0]=1;ram[3][1]=1;ram[3][2]=0;ram[3][3]=1;ram[3][4]=1;ram[3][5]=1;ram[3][6]=1;ram[3][7]=1;ram[3][8]=1;ram[3][9]=0;ram[3][10]=1;ram[3][11]=1;ram[3][12]=1;ram[3][13]=0;ram[3][14]=0;ram[3][15]=0;ram[3][16]=1;ram[3][17]=1;ram[3][18]=0;ram[3][19]=1;ram[3][20]=1;ram[3][21]=1;ram[3][22]=0;ram[3][23]=0;ram[3][24]=1;ram[3][25]=1;ram[3][26]=1;ram[3][27]=0;ram[3][28]=0;ram[3][29]=0;ram[3][30]=0;ram[3][31]=1;ram[3][32]=0;ram[3][33]=1;ram[3][34]=1;ram[3][35]=1;ram[3][36]=1;ram[3][37]=1;ram[3][38]=1;ram[3][39]=0;ram[3][40]=1;ram[3][41]=1;ram[3][42]=1;ram[3][43]=0;ram[3][44]=1;ram[3][45]=0;ram[3][46]=0;ram[3][47]=1;ram[3][48]=0;ram[3][49]=0;ram[3][50]=1;ram[3][51]=1;ram[3][52]=1;ram[3][53]=0;ram[3][54]=1;ram[3][55]=1;ram[3][56]=0;ram[3][57]=0;ram[3][58]=0;ram[3][59]=0;ram[3][60]=1;ram[3][61]=0;ram[3][62]=0;ram[3][63]=0;ram[3][64]=1;ram[3][65]=1;ram[3][66]=1;ram[3][67]=0;ram[3][68]=1;ram[3][69]=1;ram[3][70]=0;ram[3][71]=0;ram[3][72]=1;ram[3][73]=0;ram[3][74]=1;ram[3][75]=1;ram[3][76]=1;ram[3][77]=1;ram[3][78]=0;ram[3][79]=0;ram[3][80]=1;ram[3][81]=1;ram[3][82]=1;ram[3][83]=0;ram[3][84]=0;ram[3][85]=0;ram[3][86]=1;ram[3][87]=1;ram[3][88]=0;ram[3][89]=1;ram[3][90]=0;ram[3][91]=0;ram[3][92]=1;ram[3][93]=1;ram[3][94]=0;ram[3][95]=1;ram[3][96]=1;ram[3][97]=1;ram[3][98]=0;ram[3][99]=0;ram[3][100]=0;ram[3][101]=1;ram[3][102]=0;ram[3][103]=1;ram[3][104]=1;ram[3][105]=0;ram[3][106]=1;ram[3][107]=1;ram[3][108]=0;ram[3][109]=1;ram[3][110]=1;ram[3][111]=0;ram[3][112]=0;ram[3][113]=1;ram[3][114]=1;ram[3][115]=0;ram[3][116]=1;ram[3][117]=1;ram[3][118]=1;ram[3][119]=1;ram[3][120]=1;ram[3][121]=1;ram[3][122]=0;ram[3][123]=1;ram[3][124]=1;ram[3][125]=0;ram[3][126]=0;ram[3][127]=1;ram[3][128]=0;ram[3][129]=1;ram[3][130]=1;ram[3][131]=0;ram[3][132]=1;ram[3][133]=1;ram[3][134]=1;ram[3][135]=0;ram[3][136]=0;
        ram[4][0]=1;ram[4][1]=1;ram[4][2]=1;ram[4][3]=1;ram[4][4]=1;ram[4][5]=1;ram[4][6]=0;ram[4][7]=0;ram[4][8]=0;ram[4][9]=0;ram[4][10]=1;ram[4][11]=0;ram[4][12]=1;ram[4][13]=1;ram[4][14]=1;ram[4][15]=0;ram[4][16]=1;ram[4][17]=0;ram[4][18]=1;ram[4][19]=1;ram[4][20]=1;ram[4][21]=1;ram[4][22]=0;ram[4][23]=1;ram[4][24]=0;ram[4][25]=1;ram[4][26]=1;ram[4][27]=1;ram[4][28]=1;ram[4][29]=0;ram[4][30]=0;ram[4][31]=1;ram[4][32]=1;ram[4][33]=1;ram[4][34]=1;ram[4][35]=0;ram[4][36]=1;ram[4][37]=1;ram[4][38]=0;ram[4][39]=0;ram[4][40]=0;ram[4][41]=1;ram[4][42]=0;ram[4][43]=1;ram[4][44]=1;ram[4][45]=1;ram[4][46]=0;ram[4][47]=1;ram[4][48]=1;ram[4][49]=0;ram[4][50]=0;ram[4][51]=1;ram[4][52]=1;ram[4][53]=1;ram[4][54]=1;ram[4][55]=1;ram[4][56]=1;ram[4][57]=1;ram[4][58]=1;ram[4][59]=0;ram[4][60]=1;ram[4][61]=1;ram[4][62]=0;ram[4][63]=1;ram[4][64]=1;ram[4][65]=1;ram[4][66]=1;ram[4][67]=1;ram[4][68]=0;ram[4][69]=0;ram[4][70]=0;ram[4][71]=1;ram[4][72]=0;ram[4][73]=0;ram[4][74]=0;ram[4][75]=1;ram[4][76]=1;ram[4][77]=1;ram[4][78]=1;ram[4][79]=1;ram[4][80]=1;ram[4][81]=1;ram[4][82]=0;ram[4][83]=1;ram[4][84]=1;ram[4][85]=0;ram[4][86]=0;ram[4][87]=1;ram[4][88]=1;ram[4][89]=1;ram[4][90]=0;ram[4][91]=1;ram[4][92]=1;ram[4][93]=0;ram[4][94]=1;ram[4][95]=1;ram[4][96]=0;ram[4][97]=0;ram[4][98]=0;ram[4][99]=1;ram[4][100]=0;ram[4][101]=0;ram[4][102]=1;ram[4][103]=1;ram[4][104]=0;ram[4][105]=1;ram[4][106]=1;ram[4][107]=1;ram[4][108]=1;ram[4][109]=1;ram[4][110]=0;ram[4][111]=0;ram[4][112]=1;ram[4][113]=1;ram[4][114]=0;ram[4][115]=1;ram[4][116]=0;ram[4][117]=0;ram[4][118]=0;ram[4][119]=1;ram[4][120]=0;ram[4][121]=1;ram[4][122]=1;ram[4][123]=1;ram[4][124]=1;ram[4][125]=0;ram[4][126]=0;ram[4][127]=1;ram[4][128]=0;ram[4][129]=1;ram[4][130]=1;ram[4][131]=0;ram[4][132]=0;ram[4][133]=1;ram[4][134]=1;ram[4][135]=0;ram[4][136]=1;
        ram[5][0]=1;ram[5][1]=0;ram[5][2]=1;ram[5][3]=0;ram[5][4]=0;ram[5][5]=1;ram[5][6]=0;ram[5][7]=1;ram[5][8]=0;ram[5][9]=1;ram[5][10]=1;ram[5][11]=0;ram[5][12]=1;ram[5][13]=0;ram[5][14]=0;ram[5][15]=1;ram[5][16]=1;ram[5][17]=0;ram[5][18]=0;ram[5][19]=1;ram[5][20]=1;ram[5][21]=1;ram[5][22]=1;ram[5][23]=1;ram[5][24]=1;ram[5][25]=0;ram[5][26]=1;ram[5][27]=1;ram[5][28]=0;ram[5][29]=1;ram[5][30]=1;ram[5][31]=1;ram[5][32]=1;ram[5][33]=1;ram[5][34]=1;ram[5][35]=0;ram[5][36]=1;ram[5][37]=1;ram[5][38]=0;ram[5][39]=0;ram[5][40]=1;ram[5][41]=1;ram[5][42]=1;ram[5][43]=1;ram[5][44]=0;ram[5][45]=0;ram[5][46]=1;ram[5][47]=1;ram[5][48]=0;ram[5][49]=1;ram[5][50]=0;ram[5][51]=1;ram[5][52]=1;ram[5][53]=0;ram[5][54]=0;ram[5][55]=0;ram[5][56]=1;ram[5][57]=1;ram[5][58]=1;ram[5][59]=1;ram[5][60]=1;ram[5][61]=1;ram[5][62]=1;ram[5][63]=1;ram[5][64]=0;ram[5][65]=1;ram[5][66]=1;ram[5][67]=1;ram[5][68]=0;ram[5][69]=0;ram[5][70]=1;ram[5][71]=1;ram[5][72]=1;ram[5][73]=1;ram[5][74]=1;ram[5][75]=1;ram[5][76]=0;ram[5][77]=1;ram[5][78]=1;ram[5][79]=0;ram[5][80]=1;ram[5][81]=0;ram[5][82]=0;ram[5][83]=1;ram[5][84]=1;ram[5][85]=0;ram[5][86]=0;ram[5][87]=0;ram[5][88]=1;ram[5][89]=1;ram[5][90]=0;ram[5][91]=1;ram[5][92]=0;ram[5][93]=1;ram[5][94]=0;ram[5][95]=0;ram[5][96]=0;ram[5][97]=1;ram[5][98]=0;ram[5][99]=1;ram[5][100]=0;ram[5][101]=0;ram[5][102]=0;ram[5][103]=1;ram[5][104]=1;ram[5][105]=1;ram[5][106]=1;ram[5][107]=1;ram[5][108]=1;ram[5][109]=1;ram[5][110]=1;ram[5][111]=1;ram[5][112]=0;ram[5][113]=1;ram[5][114]=0;ram[5][115]=0;ram[5][116]=0;ram[5][117]=1;ram[5][118]=0;ram[5][119]=0;ram[5][120]=0;ram[5][121]=1;ram[5][122]=1;ram[5][123]=1;ram[5][124]=1;ram[5][125]=0;ram[5][126]=1;ram[5][127]=1;ram[5][128]=1;ram[5][129]=1;ram[5][130]=0;ram[5][131]=1;ram[5][132]=1;ram[5][133]=1;ram[5][134]=1;ram[5][135]=0;ram[5][136]=0;
        ram[6][0]=1;ram[6][1]=1;ram[6][2]=0;ram[6][3]=0;ram[6][4]=0;ram[6][5]=1;ram[6][6]=1;ram[6][7]=1;ram[6][8]=1;ram[6][9]=1;ram[6][10]=1;ram[6][11]=0;ram[6][12]=1;ram[6][13]=0;ram[6][14]=0;ram[6][15]=1;ram[6][16]=0;ram[6][17]=1;ram[6][18]=1;ram[6][19]=0;ram[6][20]=0;ram[6][21]=1;ram[6][22]=1;ram[6][23]=0;ram[6][24]=0;ram[6][25]=1;ram[6][26]=0;ram[6][27]=1;ram[6][28]=0;ram[6][29]=1;ram[6][30]=1;ram[6][31]=1;ram[6][32]=0;ram[6][33]=0;ram[6][34]=1;ram[6][35]=0;ram[6][36]=1;ram[6][37]=0;ram[6][38]=1;ram[6][39]=1;ram[6][40]=1;ram[6][41]=1;ram[6][42]=0;ram[6][43]=1;ram[6][44]=1;ram[6][45]=1;ram[6][46]=0;ram[6][47]=1;ram[6][48]=1;ram[6][49]=1;ram[6][50]=1;ram[6][51]=1;ram[6][52]=1;ram[6][53]=1;ram[6][54]=0;ram[6][55]=0;ram[6][56]=0;ram[6][57]=1;ram[6][58]=0;ram[6][59]=1;ram[6][60]=0;ram[6][61]=1;ram[6][62]=1;ram[6][63]=1;ram[6][64]=1;ram[6][65]=1;ram[6][66]=1;ram[6][67]=0;ram[6][68]=1;ram[6][69]=1;ram[6][70]=1;ram[6][71]=0;ram[6][72]=0;ram[6][73]=0;ram[6][74]=1;ram[6][75]=1;ram[6][76]=1;ram[6][77]=1;ram[6][78]=1;ram[6][79]=0;ram[6][80]=1;ram[6][81]=1;ram[6][82]=0;ram[6][83]=0;ram[6][84]=1;ram[6][85]=0;ram[6][86]=0;ram[6][87]=1;ram[6][88]=1;ram[6][89]=1;ram[6][90]=1;ram[6][91]=0;ram[6][92]=1;ram[6][93]=1;ram[6][94]=0;ram[6][95]=0;ram[6][96]=1;ram[6][97]=1;ram[6][98]=1;ram[6][99]=1;ram[6][100]=1;ram[6][101]=1;ram[6][102]=1;ram[6][103]=1;ram[6][104]=0;ram[6][105]=0;ram[6][106]=0;ram[6][107]=1;ram[6][108]=0;ram[6][109]=1;ram[6][110]=0;ram[6][111]=1;ram[6][112]=0;ram[6][113]=0;ram[6][114]=0;ram[6][115]=1;ram[6][116]=1;ram[6][117]=1;ram[6][118]=1;ram[6][119]=0;ram[6][120]=0;ram[6][121]=1;ram[6][122]=1;ram[6][123]=0;ram[6][124]=1;ram[6][125]=1;ram[6][126]=1;ram[6][127]=1;ram[6][128]=0;ram[6][129]=1;ram[6][130]=1;ram[6][131]=1;ram[6][132]=1;ram[6][133]=1;ram[6][134]=1;ram[6][135]=1;ram[6][136]=1;
        ram[7][0]=1;ram[7][1]=1;ram[7][2]=1;ram[7][3]=1;ram[7][4]=0;ram[7][5]=1;ram[7][6]=1;ram[7][7]=1;ram[7][8]=1;ram[7][9]=0;ram[7][10]=1;ram[7][11]=1;ram[7][12]=0;ram[7][13]=1;ram[7][14]=0;ram[7][15]=1;ram[7][16]=1;ram[7][17]=1;ram[7][18]=1;ram[7][19]=1;ram[7][20]=1;ram[7][21]=1;ram[7][22]=1;ram[7][23]=0;ram[7][24]=0;ram[7][25]=1;ram[7][26]=0;ram[7][27]=0;ram[7][28]=1;ram[7][29]=1;ram[7][30]=1;ram[7][31]=1;ram[7][32]=0;ram[7][33]=0;ram[7][34]=0;ram[7][35]=1;ram[7][36]=1;ram[7][37]=1;ram[7][38]=1;ram[7][39]=1;ram[7][40]=0;ram[7][41]=0;ram[7][42]=1;ram[7][43]=1;ram[7][44]=1;ram[7][45]=1;ram[7][46]=0;ram[7][47]=1;ram[7][48]=0;ram[7][49]=0;ram[7][50]=1;ram[7][51]=0;ram[7][52]=0;ram[7][53]=0;ram[7][54]=0;ram[7][55]=1;ram[7][56]=1;ram[7][57]=1;ram[7][58]=1;ram[7][59]=1;ram[7][60]=1;ram[7][61]=1;ram[7][62]=1;ram[7][63]=0;ram[7][64]=1;ram[7][65]=0;ram[7][66]=1;ram[7][67]=0;ram[7][68]=0;ram[7][69]=1;ram[7][70]=1;ram[7][71]=0;ram[7][72]=0;ram[7][73]=0;ram[7][74]=1;ram[7][75]=1;ram[7][76]=0;ram[7][77]=0;ram[7][78]=1;ram[7][79]=1;ram[7][80]=1;ram[7][81]=1;ram[7][82]=1;ram[7][83]=0;ram[7][84]=1;ram[7][85]=0;ram[7][86]=1;ram[7][87]=0;ram[7][88]=0;ram[7][89]=0;ram[7][90]=1;ram[7][91]=1;ram[7][92]=1;ram[7][93]=0;ram[7][94]=1;ram[7][95]=1;ram[7][96]=1;ram[7][97]=1;ram[7][98]=1;ram[7][99]=1;ram[7][100]=1;ram[7][101]=1;ram[7][102]=1;ram[7][103]=1;ram[7][104]=1;ram[7][105]=0;ram[7][106]=1;ram[7][107]=0;ram[7][108]=1;ram[7][109]=0;ram[7][110]=0;ram[7][111]=1;ram[7][112]=0;ram[7][113]=1;ram[7][114]=1;ram[7][115]=1;ram[7][116]=0;ram[7][117]=0;ram[7][118]=1;ram[7][119]=1;ram[7][120]=0;ram[7][121]=1;ram[7][122]=1;ram[7][123]=0;ram[7][124]=0;ram[7][125]=1;ram[7][126]=1;ram[7][127]=1;ram[7][128]=1;ram[7][129]=1;ram[7][130]=1;ram[7][131]=1;ram[7][132]=1;ram[7][133]=0;ram[7][134]=0;ram[7][135]=1;ram[7][136]=0;
        ram[8][0]=1;ram[8][1]=1;ram[8][2]=0;ram[8][3]=1;ram[8][4]=0;ram[8][5]=0;ram[8][6]=1;ram[8][7]=1;ram[8][8]=0;ram[8][9]=1;ram[8][10]=1;ram[8][11]=1;ram[8][12]=1;ram[8][13]=1;ram[8][14]=1;ram[8][15]=0;ram[8][16]=0;ram[8][17]=1;ram[8][18]=0;ram[8][19]=1;ram[8][20]=1;ram[8][21]=1;ram[8][22]=1;ram[8][23]=1;ram[8][24]=1;ram[8][25]=0;ram[8][26]=0;ram[8][27]=1;ram[8][28]=1;ram[8][29]=0;ram[8][30]=1;ram[8][31]=1;ram[8][32]=0;ram[8][33]=1;ram[8][34]=1;ram[8][35]=1;ram[8][36]=0;ram[8][37]=1;ram[8][38]=0;ram[8][39]=1;ram[8][40]=0;ram[8][41]=1;ram[8][42]=1;ram[8][43]=0;ram[8][44]=0;ram[8][45]=1;ram[8][46]=1;ram[8][47]=1;ram[8][48]=0;ram[8][49]=1;ram[8][50]=0;ram[8][51]=1;ram[8][52]=1;ram[8][53]=1;ram[8][54]=1;ram[8][55]=1;ram[8][56]=1;ram[8][57]=0;ram[8][58]=1;ram[8][59]=1;ram[8][60]=1;ram[8][61]=1;ram[8][62]=0;ram[8][63]=0;ram[8][64]=1;ram[8][65]=1;ram[8][66]=1;ram[8][67]=1;ram[8][68]=1;ram[8][69]=1;ram[8][70]=1;ram[8][71]=1;ram[8][72]=1;ram[8][73]=1;ram[8][74]=1;ram[8][75]=1;ram[8][76]=1;ram[8][77]=1;ram[8][78]=1;ram[8][79]=0;ram[8][80]=0;ram[8][81]=1;ram[8][82]=1;ram[8][83]=1;ram[8][84]=0;ram[8][85]=1;ram[8][86]=0;ram[8][87]=1;ram[8][88]=1;ram[8][89]=1;ram[8][90]=1;ram[8][91]=0;ram[8][92]=0;ram[8][93]=1;ram[8][94]=0;ram[8][95]=0;ram[8][96]=0;ram[8][97]=1;ram[8][98]=1;ram[8][99]=1;ram[8][100]=1;ram[8][101]=1;ram[8][102]=1;ram[8][103]=1;ram[8][104]=1;ram[8][105]=1;ram[8][106]=1;ram[8][107]=1;ram[8][108]=1;ram[8][109]=0;ram[8][110]=1;ram[8][111]=0;ram[8][112]=0;ram[8][113]=0;ram[8][114]=1;ram[8][115]=1;ram[8][116]=0;ram[8][117]=0;ram[8][118]=1;ram[8][119]=1;ram[8][120]=0;ram[8][121]=1;ram[8][122]=1;ram[8][123]=1;ram[8][124]=0;ram[8][125]=0;ram[8][126]=1;ram[8][127]=0;ram[8][128]=1;ram[8][129]=1;ram[8][130]=1;ram[8][131]=1;ram[8][132]=0;ram[8][133]=1;ram[8][134]=1;ram[8][135]=0;ram[8][136]=1;
        ram[9][0]=1;ram[9][1]=0;ram[9][2]=1;ram[9][3]=1;ram[9][4]=1;ram[9][5]=0;ram[9][6]=1;ram[9][7]=1;ram[9][8]=0;ram[9][9]=1;ram[9][10]=0;ram[9][11]=1;ram[9][12]=1;ram[9][13]=0;ram[9][14]=1;ram[9][15]=0;ram[9][16]=1;ram[9][17]=1;ram[9][18]=1;ram[9][19]=1;ram[9][20]=1;ram[9][21]=1;ram[9][22]=0;ram[9][23]=1;ram[9][24]=1;ram[9][25]=1;ram[9][26]=1;ram[9][27]=0;ram[9][28]=1;ram[9][29]=0;ram[9][30]=0;ram[9][31]=0;ram[9][32]=0;ram[9][33]=1;ram[9][34]=1;ram[9][35]=1;ram[9][36]=0;ram[9][37]=1;ram[9][38]=1;ram[9][39]=0;ram[9][40]=1;ram[9][41]=1;ram[9][42]=1;ram[9][43]=1;ram[9][44]=1;ram[9][45]=0;ram[9][46]=1;ram[9][47]=1;ram[9][48]=1;ram[9][49]=0;ram[9][50]=1;ram[9][51]=0;ram[9][52]=1;ram[9][53]=1;ram[9][54]=0;ram[9][55]=0;ram[9][56]=0;ram[9][57]=1;ram[9][58]=1;ram[9][59]=0;ram[9][60]=1;ram[9][61]=1;ram[9][62]=1;ram[9][63]=0;ram[9][64]=1;ram[9][65]=1;ram[9][66]=1;ram[9][67]=1;ram[9][68]=1;ram[9][69]=0;ram[9][70]=1;ram[9][71]=1;ram[9][72]=1;ram[9][73]=1;ram[9][74]=0;ram[9][75]=1;ram[9][76]=0;ram[9][77]=1;ram[9][78]=0;ram[9][79]=1;ram[9][80]=1;ram[9][81]=1;ram[9][82]=1;ram[9][83]=1;ram[9][84]=0;ram[9][85]=0;ram[9][86]=0;ram[9][87]=1;ram[9][88]=1;ram[9][89]=0;ram[9][90]=0;ram[9][91]=0;ram[9][92]=1;ram[9][93]=1;ram[9][94]=0;ram[9][95]=1;ram[9][96]=0;ram[9][97]=1;ram[9][98]=0;ram[9][99]=1;ram[9][100]=0;ram[9][101]=1;ram[9][102]=1;ram[9][103]=1;ram[9][104]=1;ram[9][105]=1;ram[9][106]=0;ram[9][107]=1;ram[9][108]=1;ram[9][109]=1;ram[9][110]=1;ram[9][111]=0;ram[9][112]=1;ram[9][113]=1;ram[9][114]=1;ram[9][115]=0;ram[9][116]=1;ram[9][117]=1;ram[9][118]=1;ram[9][119]=0;ram[9][120]=0;ram[9][121]=1;ram[9][122]=0;ram[9][123]=0;ram[9][124]=0;ram[9][125]=1;ram[9][126]=1;ram[9][127]=1;ram[9][128]=1;ram[9][129]=1;ram[9][130]=1;ram[9][131]=0;ram[9][132]=1;ram[9][133]=0;ram[9][134]=1;ram[9][135]=1;ram[9][136]=1;
        ram[10][0]=1;ram[10][1]=1;ram[10][2]=1;ram[10][3]=1;ram[10][4]=0;ram[10][5]=1;ram[10][6]=1;ram[10][7]=1;ram[10][8]=1;ram[10][9]=1;ram[10][10]=1;ram[10][11]=1;ram[10][12]=1;ram[10][13]=1;ram[10][14]=1;ram[10][15]=1;ram[10][16]=1;ram[10][17]=0;ram[10][18]=1;ram[10][19]=1;ram[10][20]=1;ram[10][21]=1;ram[10][22]=1;ram[10][23]=1;ram[10][24]=1;ram[10][25]=1;ram[10][26]=0;ram[10][27]=0;ram[10][28]=0;ram[10][29]=1;ram[10][30]=1;ram[10][31]=1;ram[10][32]=0;ram[10][33]=0;ram[10][34]=1;ram[10][35]=1;ram[10][36]=0;ram[10][37]=1;ram[10][38]=0;ram[10][39]=1;ram[10][40]=0;ram[10][41]=1;ram[10][42]=1;ram[10][43]=0;ram[10][44]=1;ram[10][45]=0;ram[10][46]=0;ram[10][47]=1;ram[10][48]=0;ram[10][49]=1;ram[10][50]=1;ram[10][51]=1;ram[10][52]=1;ram[10][53]=1;ram[10][54]=0;ram[10][55]=1;ram[10][56]=1;ram[10][57]=0;ram[10][58]=0;ram[10][59]=0;ram[10][60]=1;ram[10][61]=1;ram[10][62]=1;ram[10][63]=0;ram[10][64]=0;ram[10][65]=0;ram[10][66]=0;ram[10][67]=1;ram[10][68]=0;ram[10][69]=0;ram[10][70]=1;ram[10][71]=1;ram[10][72]=1;ram[10][73]=1;ram[10][74]=1;ram[10][75]=1;ram[10][76]=1;ram[10][77]=1;ram[10][78]=1;ram[10][79]=0;ram[10][80]=1;ram[10][81]=0;ram[10][82]=1;ram[10][83]=1;ram[10][84]=1;ram[10][85]=0;ram[10][86]=1;ram[10][87]=0;ram[10][88]=1;ram[10][89]=0;ram[10][90]=0;ram[10][91]=1;ram[10][92]=0;ram[10][93]=1;ram[10][94]=0;ram[10][95]=1;ram[10][96]=1;ram[10][97]=0;ram[10][98]=1;ram[10][99]=1;ram[10][100]=1;ram[10][101]=1;ram[10][102]=0;ram[10][103]=0;ram[10][104]=1;ram[10][105]=1;ram[10][106]=0;ram[10][107]=0;ram[10][108]=0;ram[10][109]=0;ram[10][110]=1;ram[10][111]=1;ram[10][112]=1;ram[10][113]=1;ram[10][114]=1;ram[10][115]=1;ram[10][116]=1;ram[10][117]=0;ram[10][118]=1;ram[10][119]=1;ram[10][120]=1;ram[10][121]=1;ram[10][122]=1;ram[10][123]=1;ram[10][124]=0;ram[10][125]=1;ram[10][126]=0;ram[10][127]=1;ram[10][128]=1;ram[10][129]=1;ram[10][130]=1;ram[10][131]=1;ram[10][132]=1;ram[10][133]=1;ram[10][134]=1;ram[10][135]=1;ram[10][136]=0;
        ram[11][0]=1;ram[11][1]=1;ram[11][2]=1;ram[11][3]=1;ram[11][4]=1;ram[11][5]=1;ram[11][6]=1;ram[11][7]=0;ram[11][8]=1;ram[11][9]=0;ram[11][10]=1;ram[11][11]=1;ram[11][12]=1;ram[11][13]=1;ram[11][14]=1;ram[11][15]=1;ram[11][16]=0;ram[11][17]=1;ram[11][18]=1;ram[11][19]=0;ram[11][20]=1;ram[11][21]=1;ram[11][22]=1;ram[11][23]=1;ram[11][24]=0;ram[11][25]=1;ram[11][26]=0;ram[11][27]=1;ram[11][28]=0;ram[11][29]=0;ram[11][30]=0;ram[11][31]=0;ram[11][32]=1;ram[11][33]=1;ram[11][34]=1;ram[11][35]=1;ram[11][36]=0;ram[11][37]=0;ram[11][38]=1;ram[11][39]=1;ram[11][40]=0;ram[11][41]=1;ram[11][42]=1;ram[11][43]=1;ram[11][44]=0;ram[11][45]=1;ram[11][46]=0;ram[11][47]=1;ram[11][48]=1;ram[11][49]=1;ram[11][50]=1;ram[11][51]=1;ram[11][52]=0;ram[11][53]=0;ram[11][54]=0;ram[11][55]=1;ram[11][56]=1;ram[11][57]=1;ram[11][58]=1;ram[11][59]=1;ram[11][60]=1;ram[11][61]=0;ram[11][62]=1;ram[11][63]=0;ram[11][64]=1;ram[11][65]=1;ram[11][66]=1;ram[11][67]=1;ram[11][68]=1;ram[11][69]=1;ram[11][70]=1;ram[11][71]=1;ram[11][72]=1;ram[11][73]=0;ram[11][74]=0;ram[11][75]=1;ram[11][76]=1;ram[11][77]=0;ram[11][78]=0;ram[11][79]=1;ram[11][80]=1;ram[11][81]=0;ram[11][82]=0;ram[11][83]=1;ram[11][84]=1;ram[11][85]=1;ram[11][86]=1;ram[11][87]=0;ram[11][88]=1;ram[11][89]=0;ram[11][90]=0;ram[11][91]=1;ram[11][92]=0;ram[11][93]=0;ram[11][94]=0;ram[11][95]=1;ram[11][96]=1;ram[11][97]=1;ram[11][98]=1;ram[11][99]=0;ram[11][100]=0;ram[11][101]=0;ram[11][102]=0;ram[11][103]=0;ram[11][104]=1;ram[11][105]=0;ram[11][106]=1;ram[11][107]=1;ram[11][108]=1;ram[11][109]=0;ram[11][110]=1;ram[11][111]=0;ram[11][112]=1;ram[11][113]=1;ram[11][114]=1;ram[11][115]=0;ram[11][116]=1;ram[11][117]=1;ram[11][118]=1;ram[11][119]=1;ram[11][120]=1;ram[11][121]=0;ram[11][122]=1;ram[11][123]=1;ram[11][124]=0;ram[11][125]=0;ram[11][126]=1;ram[11][127]=0;ram[11][128]=1;ram[11][129]=0;ram[11][130]=0;ram[11][131]=0;ram[11][132]=1;ram[11][133]=0;ram[11][134]=0;ram[11][135]=0;ram[11][136]=1;
        ram[12][0]=0;ram[12][1]=0;ram[12][2]=1;ram[12][3]=1;ram[12][4]=0;ram[12][5]=0;ram[12][6]=1;ram[12][7]=0;ram[12][8]=1;ram[12][9]=0;ram[12][10]=0;ram[12][11]=0;ram[12][12]=0;ram[12][13]=1;ram[12][14]=1;ram[12][15]=0;ram[12][16]=1;ram[12][17]=1;ram[12][18]=1;ram[12][19]=0;ram[12][20]=0;ram[12][21]=1;ram[12][22]=1;ram[12][23]=1;ram[12][24]=1;ram[12][25]=1;ram[12][26]=0;ram[12][27]=1;ram[12][28]=1;ram[12][29]=1;ram[12][30]=1;ram[12][31]=0;ram[12][32]=0;ram[12][33]=1;ram[12][34]=1;ram[12][35]=1;ram[12][36]=1;ram[12][37]=0;ram[12][38]=1;ram[12][39]=0;ram[12][40]=1;ram[12][41]=0;ram[12][42]=1;ram[12][43]=1;ram[12][44]=1;ram[12][45]=0;ram[12][46]=0;ram[12][47]=0;ram[12][48]=1;ram[12][49]=1;ram[12][50]=1;ram[12][51]=0;ram[12][52]=1;ram[12][53]=1;ram[12][54]=0;ram[12][55]=1;ram[12][56]=0;ram[12][57]=1;ram[12][58]=1;ram[12][59]=1;ram[12][60]=0;ram[12][61]=0;ram[12][62]=0;ram[12][63]=1;ram[12][64]=1;ram[12][65]=1;ram[12][66]=1;ram[12][67]=1;ram[12][68]=0;ram[12][69]=0;ram[12][70]=1;ram[12][71]=0;ram[12][72]=1;ram[12][73]=0;ram[12][74]=0;ram[12][75]=0;ram[12][76]=0;ram[12][77]=0;ram[12][78]=0;ram[12][79]=0;ram[12][80]=1;ram[12][81]=1;ram[12][82]=0;ram[12][83]=0;ram[12][84]=1;ram[12][85]=1;ram[12][86]=0;ram[12][87]=1;ram[12][88]=0;ram[12][89]=1;ram[12][90]=1;ram[12][91]=1;ram[12][92]=1;ram[12][93]=1;ram[12][94]=1;ram[12][95]=0;ram[12][96]=1;ram[12][97]=1;ram[12][98]=1;ram[12][99]=1;ram[12][100]=1;ram[12][101]=1;ram[12][102]=1;ram[12][103]=0;ram[12][104]=1;ram[12][105]=1;ram[12][106]=0;ram[12][107]=1;ram[12][108]=1;ram[12][109]=0;ram[12][110]=1;ram[12][111]=0;ram[12][112]=0;ram[12][113]=1;ram[12][114]=1;ram[12][115]=1;ram[12][116]=0;ram[12][117]=1;ram[12][118]=1;ram[12][119]=1;ram[12][120]=0;ram[12][121]=1;ram[12][122]=1;ram[12][123]=1;ram[12][124]=0;ram[12][125]=0;ram[12][126]=0;ram[12][127]=1;ram[12][128]=1;ram[12][129]=0;ram[12][130]=1;ram[12][131]=0;ram[12][132]=1;ram[12][133]=1;ram[12][134]=1;ram[12][135]=0;ram[12][136]=0;
        ram[13][0]=1;ram[13][1]=0;ram[13][2]=0;ram[13][3]=0;ram[13][4]=1;ram[13][5]=1;ram[13][6]=0;ram[13][7]=1;ram[13][8]=1;ram[13][9]=0;ram[13][10]=1;ram[13][11]=0;ram[13][12]=0;ram[13][13]=1;ram[13][14]=1;ram[13][15]=1;ram[13][16]=1;ram[13][17]=1;ram[13][18]=0;ram[13][19]=0;ram[13][20]=1;ram[13][21]=1;ram[13][22]=1;ram[13][23]=0;ram[13][24]=1;ram[13][25]=1;ram[13][26]=0;ram[13][27]=1;ram[13][28]=1;ram[13][29]=1;ram[13][30]=1;ram[13][31]=1;ram[13][32]=1;ram[13][33]=1;ram[13][34]=1;ram[13][35]=1;ram[13][36]=0;ram[13][37]=0;ram[13][38]=1;ram[13][39]=1;ram[13][40]=0;ram[13][41]=1;ram[13][42]=1;ram[13][43]=1;ram[13][44]=1;ram[13][45]=0;ram[13][46]=0;ram[13][47]=1;ram[13][48]=1;ram[13][49]=0;ram[13][50]=1;ram[13][51]=1;ram[13][52]=0;ram[13][53]=0;ram[13][54]=1;ram[13][55]=1;ram[13][56]=1;ram[13][57]=1;ram[13][58]=1;ram[13][59]=0;ram[13][60]=1;ram[13][61]=1;ram[13][62]=1;ram[13][63]=1;ram[13][64]=1;ram[13][65]=1;ram[13][66]=1;ram[13][67]=1;ram[13][68]=1;ram[13][69]=1;ram[13][70]=1;ram[13][71]=0;ram[13][72]=1;ram[13][73]=0;ram[13][74]=1;ram[13][75]=0;ram[13][76]=1;ram[13][77]=1;ram[13][78]=0;ram[13][79]=0;ram[13][80]=1;ram[13][81]=1;ram[13][82]=0;ram[13][83]=0;ram[13][84]=1;ram[13][85]=1;ram[13][86]=1;ram[13][87]=0;ram[13][88]=1;ram[13][89]=1;ram[13][90]=1;ram[13][91]=1;ram[13][92]=0;ram[13][93]=0;ram[13][94]=1;ram[13][95]=1;ram[13][96]=1;ram[13][97]=1;ram[13][98]=0;ram[13][99]=1;ram[13][100]=1;ram[13][101]=1;ram[13][102]=1;ram[13][103]=0;ram[13][104]=0;ram[13][105]=1;ram[13][106]=0;ram[13][107]=1;ram[13][108]=0;ram[13][109]=0;ram[13][110]=1;ram[13][111]=1;ram[13][112]=1;ram[13][113]=1;ram[13][114]=0;ram[13][115]=0;ram[13][116]=1;ram[13][117]=1;ram[13][118]=1;ram[13][119]=0;ram[13][120]=1;ram[13][121]=0;ram[13][122]=0;ram[13][123]=1;ram[13][124]=1;ram[13][125]=0;ram[13][126]=1;ram[13][127]=0;ram[13][128]=0;ram[13][129]=1;ram[13][130]=1;ram[13][131]=0;ram[13][132]=1;ram[13][133]=0;ram[13][134]=1;ram[13][135]=0;ram[13][136]=0;
        ram[14][0]=1;ram[14][1]=0;ram[14][2]=1;ram[14][3]=1;ram[14][4]=1;ram[14][5]=1;ram[14][6]=0;ram[14][7]=1;ram[14][8]=0;ram[14][9]=0;ram[14][10]=1;ram[14][11]=1;ram[14][12]=1;ram[14][13]=1;ram[14][14]=1;ram[14][15]=1;ram[14][16]=0;ram[14][17]=1;ram[14][18]=0;ram[14][19]=1;ram[14][20]=1;ram[14][21]=1;ram[14][22]=1;ram[14][23]=1;ram[14][24]=1;ram[14][25]=1;ram[14][26]=1;ram[14][27]=0;ram[14][28]=0;ram[14][29]=0;ram[14][30]=1;ram[14][31]=1;ram[14][32]=1;ram[14][33]=1;ram[14][34]=1;ram[14][35]=1;ram[14][36]=0;ram[14][37]=1;ram[14][38]=1;ram[14][39]=1;ram[14][40]=1;ram[14][41]=1;ram[14][42]=1;ram[14][43]=1;ram[14][44]=1;ram[14][45]=1;ram[14][46]=1;ram[14][47]=1;ram[14][48]=1;ram[14][49]=1;ram[14][50]=1;ram[14][51]=1;ram[14][52]=0;ram[14][53]=1;ram[14][54]=0;ram[14][55]=0;ram[14][56]=0;ram[14][57]=1;ram[14][58]=1;ram[14][59]=1;ram[14][60]=0;ram[14][61]=1;ram[14][62]=0;ram[14][63]=1;ram[14][64]=1;ram[14][65]=1;ram[14][66]=1;ram[14][67]=1;ram[14][68]=1;ram[14][69]=1;ram[14][70]=1;ram[14][71]=1;ram[14][72]=0;ram[14][73]=1;ram[14][74]=1;ram[14][75]=0;ram[14][76]=1;ram[14][77]=1;ram[14][78]=1;ram[14][79]=0;ram[14][80]=0;ram[14][81]=1;ram[14][82]=1;ram[14][83]=1;ram[14][84]=1;ram[14][85]=1;ram[14][86]=1;ram[14][87]=1;ram[14][88]=1;ram[14][89]=0;ram[14][90]=0;ram[14][91]=0;ram[14][92]=0;ram[14][93]=0;ram[14][94]=0;ram[14][95]=1;ram[14][96]=1;ram[14][97]=1;ram[14][98]=1;ram[14][99]=0;ram[14][100]=0;ram[14][101]=1;ram[14][102]=1;ram[14][103]=1;ram[14][104]=1;ram[14][105]=0;ram[14][106]=1;ram[14][107]=1;ram[14][108]=1;ram[14][109]=1;ram[14][110]=1;ram[14][111]=1;ram[14][112]=1;ram[14][113]=0;ram[14][114]=1;ram[14][115]=1;ram[14][116]=1;ram[14][117]=1;ram[14][118]=1;ram[14][119]=1;ram[14][120]=1;ram[14][121]=1;ram[14][122]=1;ram[14][123]=1;ram[14][124]=1;ram[14][125]=0;ram[14][126]=0;ram[14][127]=1;ram[14][128]=0;ram[14][129]=1;ram[14][130]=1;ram[14][131]=0;ram[14][132]=0;ram[14][133]=0;ram[14][134]=1;ram[14][135]=0;ram[14][136]=1;
        ram[15][0]=1;ram[15][1]=1;ram[15][2]=0;ram[15][3]=1;ram[15][4]=1;ram[15][5]=1;ram[15][6]=1;ram[15][7]=0;ram[15][8]=1;ram[15][9]=0;ram[15][10]=1;ram[15][11]=1;ram[15][12]=1;ram[15][13]=1;ram[15][14]=1;ram[15][15]=1;ram[15][16]=0;ram[15][17]=1;ram[15][18]=0;ram[15][19]=1;ram[15][20]=0;ram[15][21]=1;ram[15][22]=0;ram[15][23]=0;ram[15][24]=1;ram[15][25]=0;ram[15][26]=0;ram[15][27]=1;ram[15][28]=1;ram[15][29]=1;ram[15][30]=1;ram[15][31]=1;ram[15][32]=1;ram[15][33]=1;ram[15][34]=1;ram[15][35]=1;ram[15][36]=0;ram[15][37]=1;ram[15][38]=1;ram[15][39]=1;ram[15][40]=1;ram[15][41]=1;ram[15][42]=1;ram[15][43]=0;ram[15][44]=1;ram[15][45]=0;ram[15][46]=1;ram[15][47]=1;ram[15][48]=0;ram[15][49]=0;ram[15][50]=1;ram[15][51]=1;ram[15][52]=0;ram[15][53]=1;ram[15][54]=1;ram[15][55]=1;ram[15][56]=1;ram[15][57]=1;ram[15][58]=0;ram[15][59]=0;ram[15][60]=1;ram[15][61]=1;ram[15][62]=1;ram[15][63]=1;ram[15][64]=1;ram[15][65]=1;ram[15][66]=1;ram[15][67]=0;ram[15][68]=0;ram[15][69]=1;ram[15][70]=1;ram[15][71]=0;ram[15][72]=1;ram[15][73]=1;ram[15][74]=1;ram[15][75]=1;ram[15][76]=1;ram[15][77]=1;ram[15][78]=0;ram[15][79]=0;ram[15][80]=0;ram[15][81]=1;ram[15][82]=1;ram[15][83]=1;ram[15][84]=0;ram[15][85]=1;ram[15][86]=1;ram[15][87]=0;ram[15][88]=1;ram[15][89]=1;ram[15][90]=1;ram[15][91]=1;ram[15][92]=0;ram[15][93]=0;ram[15][94]=1;ram[15][95]=0;ram[15][96]=1;ram[15][97]=1;ram[15][98]=0;ram[15][99]=1;ram[15][100]=0;ram[15][101]=1;ram[15][102]=1;ram[15][103]=1;ram[15][104]=0;ram[15][105]=1;ram[15][106]=1;ram[15][107]=1;ram[15][108]=1;ram[15][109]=1;ram[15][110]=1;ram[15][111]=1;ram[15][112]=0;ram[15][113]=0;ram[15][114]=1;ram[15][115]=1;ram[15][116]=1;ram[15][117]=1;ram[15][118]=0;ram[15][119]=1;ram[15][120]=0;ram[15][121]=1;ram[15][122]=1;ram[15][123]=1;ram[15][124]=1;ram[15][125]=1;ram[15][126]=1;ram[15][127]=1;ram[15][128]=1;ram[15][129]=0;ram[15][130]=0;ram[15][131]=0;ram[15][132]=1;ram[15][133]=1;ram[15][134]=1;ram[15][135]=0;ram[15][136]=0;
        ram[16][0]=1;ram[16][1]=0;ram[16][2]=1;ram[16][3]=0;ram[16][4]=1;ram[16][5]=0;ram[16][6]=0;ram[16][7]=1;ram[16][8]=1;ram[16][9]=0;ram[16][10]=0;ram[16][11]=0;ram[16][12]=1;ram[16][13]=1;ram[16][14]=1;ram[16][15]=1;ram[16][16]=0;ram[16][17]=1;ram[16][18]=0;ram[16][19]=0;ram[16][20]=1;ram[16][21]=1;ram[16][22]=1;ram[16][23]=1;ram[16][24]=0;ram[16][25]=1;ram[16][26]=1;ram[16][27]=1;ram[16][28]=0;ram[16][29]=0;ram[16][30]=1;ram[16][31]=1;ram[16][32]=1;ram[16][33]=0;ram[16][34]=1;ram[16][35]=1;ram[16][36]=1;ram[16][37]=1;ram[16][38]=0;ram[16][39]=1;ram[16][40]=1;ram[16][41]=1;ram[16][42]=1;ram[16][43]=1;ram[16][44]=0;ram[16][45]=1;ram[16][46]=1;ram[16][47]=1;ram[16][48]=1;ram[16][49]=0;ram[16][50]=1;ram[16][51]=1;ram[16][52]=1;ram[16][53]=0;ram[16][54]=0;ram[16][55]=1;ram[16][56]=1;ram[16][57]=0;ram[16][58]=1;ram[16][59]=1;ram[16][60]=0;ram[16][61]=1;ram[16][62]=1;ram[16][63]=1;ram[16][64]=1;ram[16][65]=1;ram[16][66]=0;ram[16][67]=0;ram[16][68]=1;ram[16][69]=0;ram[16][70]=1;ram[16][71]=1;ram[16][72]=0;ram[16][73]=1;ram[16][74]=1;ram[16][75]=0;ram[16][76]=0;ram[16][77]=0;ram[16][78]=0;ram[16][79]=1;ram[16][80]=1;ram[16][81]=0;ram[16][82]=1;ram[16][83]=1;ram[16][84]=0;ram[16][85]=0;ram[16][86]=1;ram[16][87]=1;ram[16][88]=0;ram[16][89]=1;ram[16][90]=0;ram[16][91]=0;ram[16][92]=1;ram[16][93]=1;ram[16][94]=0;ram[16][95]=1;ram[16][96]=1;ram[16][97]=0;ram[16][98]=1;ram[16][99]=1;ram[16][100]=1;ram[16][101]=1;ram[16][102]=1;ram[16][103]=1;ram[16][104]=0;ram[16][105]=1;ram[16][106]=1;ram[16][107]=1;ram[16][108]=1;ram[16][109]=0;ram[16][110]=1;ram[16][111]=0;ram[16][112]=0;ram[16][113]=1;ram[16][114]=1;ram[16][115]=1;ram[16][116]=0;ram[16][117]=1;ram[16][118]=0;ram[16][119]=1;ram[16][120]=0;ram[16][121]=1;ram[16][122]=1;ram[16][123]=1;ram[16][124]=1;ram[16][125]=1;ram[16][126]=1;ram[16][127]=1;ram[16][128]=1;ram[16][129]=0;ram[16][130]=0;ram[16][131]=0;ram[16][132]=0;ram[16][133]=1;ram[16][134]=1;ram[16][135]=0;ram[16][136]=0;
        ram[17][0]=1;ram[17][1]=1;ram[17][2]=1;ram[17][3]=0;ram[17][4]=1;ram[17][5]=1;ram[17][6]=0;ram[17][7]=0;ram[17][8]=1;ram[17][9]=1;ram[17][10]=1;ram[17][11]=0;ram[17][12]=1;ram[17][13]=1;ram[17][14]=1;ram[17][15]=0;ram[17][16]=0;ram[17][17]=0;ram[17][18]=1;ram[17][19]=0;ram[17][20]=1;ram[17][21]=1;ram[17][22]=1;ram[17][23]=1;ram[17][24]=1;ram[17][25]=1;ram[17][26]=1;ram[17][27]=0;ram[17][28]=1;ram[17][29]=0;ram[17][30]=0;ram[17][31]=1;ram[17][32]=1;ram[17][33]=1;ram[17][34]=1;ram[17][35]=1;ram[17][36]=0;ram[17][37]=1;ram[17][38]=1;ram[17][39]=1;ram[17][40]=1;ram[17][41]=0;ram[17][42]=0;ram[17][43]=0;ram[17][44]=1;ram[17][45]=0;ram[17][46]=0;ram[17][47]=0;ram[17][48]=1;ram[17][49]=1;ram[17][50]=1;ram[17][51]=0;ram[17][52]=1;ram[17][53]=0;ram[17][54]=0;ram[17][55]=1;ram[17][56]=1;ram[17][57]=1;ram[17][58]=0;ram[17][59]=0;ram[17][60]=1;ram[17][61]=0;ram[17][62]=1;ram[17][63]=0;ram[17][64]=1;ram[17][65]=0;ram[17][66]=1;ram[17][67]=1;ram[17][68]=1;ram[17][69]=0;ram[17][70]=0;ram[17][71]=1;ram[17][72]=1;ram[17][73]=1;ram[17][74]=1;ram[17][75]=1;ram[17][76]=1;ram[17][77]=1;ram[17][78]=1;ram[17][79]=0;ram[17][80]=1;ram[17][81]=1;ram[17][82]=0;ram[17][83]=1;ram[17][84]=0;ram[17][85]=1;ram[17][86]=0;ram[17][87]=1;ram[17][88]=0;ram[17][89]=0;ram[17][90]=1;ram[17][91]=0;ram[17][92]=1;ram[17][93]=1;ram[17][94]=1;ram[17][95]=1;ram[17][96]=0;ram[17][97]=1;ram[17][98]=0;ram[17][99]=1;ram[17][100]=0;ram[17][101]=1;ram[17][102]=1;ram[17][103]=1;ram[17][104]=1;ram[17][105]=1;ram[17][106]=1;ram[17][107]=1;ram[17][108]=1;ram[17][109]=1;ram[17][110]=1;ram[17][111]=0;ram[17][112]=1;ram[17][113]=1;ram[17][114]=0;ram[17][115]=1;ram[17][116]=1;ram[17][117]=1;ram[17][118]=1;ram[17][119]=0;ram[17][120]=1;ram[17][121]=1;ram[17][122]=1;ram[17][123]=0;ram[17][124]=1;ram[17][125]=1;ram[17][126]=1;ram[17][127]=1;ram[17][128]=1;ram[17][129]=1;ram[17][130]=1;ram[17][131]=1;ram[17][132]=1;ram[17][133]=0;ram[17][134]=1;ram[17][135]=0;ram[17][136]=1;
        ram[18][0]=1;ram[18][1]=1;ram[18][2]=0;ram[18][3]=1;ram[18][4]=0;ram[18][5]=0;ram[18][6]=1;ram[18][7]=1;ram[18][8]=1;ram[18][9]=1;ram[18][10]=1;ram[18][11]=1;ram[18][12]=1;ram[18][13]=1;ram[18][14]=0;ram[18][15]=1;ram[18][16]=1;ram[18][17]=1;ram[18][18]=0;ram[18][19]=1;ram[18][20]=0;ram[18][21]=1;ram[18][22]=1;ram[18][23]=0;ram[18][24]=1;ram[18][25]=1;ram[18][26]=0;ram[18][27]=0;ram[18][28]=1;ram[18][29]=1;ram[18][30]=0;ram[18][31]=1;ram[18][32]=1;ram[18][33]=0;ram[18][34]=0;ram[18][35]=1;ram[18][36]=1;ram[18][37]=1;ram[18][38]=1;ram[18][39]=0;ram[18][40]=1;ram[18][41]=1;ram[18][42]=0;ram[18][43]=1;ram[18][44]=1;ram[18][45]=1;ram[18][46]=1;ram[18][47]=1;ram[18][48]=0;ram[18][49]=1;ram[18][50]=0;ram[18][51]=0;ram[18][52]=1;ram[18][53]=0;ram[18][54]=0;ram[18][55]=1;ram[18][56]=1;ram[18][57]=1;ram[18][58]=1;ram[18][59]=1;ram[18][60]=1;ram[18][61]=1;ram[18][62]=0;ram[18][63]=0;ram[18][64]=1;ram[18][65]=0;ram[18][66]=0;ram[18][67]=1;ram[18][68]=1;ram[18][69]=1;ram[18][70]=0;ram[18][71]=0;ram[18][72]=1;ram[18][73]=0;ram[18][74]=1;ram[18][75]=0;ram[18][76]=0;ram[18][77]=1;ram[18][78]=1;ram[18][79]=0;ram[18][80]=1;ram[18][81]=1;ram[18][82]=0;ram[18][83]=1;ram[18][84]=1;ram[18][85]=1;ram[18][86]=1;ram[18][87]=0;ram[18][88]=0;ram[18][89]=1;ram[18][90]=1;ram[18][91]=1;ram[18][92]=0;ram[18][93]=0;ram[18][94]=1;ram[18][95]=1;ram[18][96]=1;ram[18][97]=0;ram[18][98]=1;ram[18][99]=1;ram[18][100]=0;ram[18][101]=1;ram[18][102]=0;ram[18][103]=1;ram[18][104]=1;ram[18][105]=1;ram[18][106]=1;ram[18][107]=1;ram[18][108]=1;ram[18][109]=0;ram[18][110]=0;ram[18][111]=0;ram[18][112]=0;ram[18][113]=1;ram[18][114]=0;ram[18][115]=0;ram[18][116]=1;ram[18][117]=1;ram[18][118]=1;ram[18][119]=0;ram[18][120]=1;ram[18][121]=1;ram[18][122]=0;ram[18][123]=1;ram[18][124]=0;ram[18][125]=0;ram[18][126]=1;ram[18][127]=0;ram[18][128]=0;ram[18][129]=1;ram[18][130]=1;ram[18][131]=1;ram[18][132]=1;ram[18][133]=0;ram[18][134]=1;ram[18][135]=0;ram[18][136]=1;
        ram[19][0]=1;ram[19][1]=0;ram[19][2]=1;ram[19][3]=0;ram[19][4]=0;ram[19][5]=1;ram[19][6]=1;ram[19][7]=1;ram[19][8]=0;ram[19][9]=0;ram[19][10]=1;ram[19][11]=1;ram[19][12]=1;ram[19][13]=1;ram[19][14]=1;ram[19][15]=1;ram[19][16]=0;ram[19][17]=0;ram[19][18]=1;ram[19][19]=1;ram[19][20]=1;ram[19][21]=0;ram[19][22]=1;ram[19][23]=1;ram[19][24]=1;ram[19][25]=1;ram[19][26]=0;ram[19][27]=1;ram[19][28]=0;ram[19][29]=0;ram[19][30]=1;ram[19][31]=1;ram[19][32]=1;ram[19][33]=0;ram[19][34]=1;ram[19][35]=0;ram[19][36]=1;ram[19][37]=0;ram[19][38]=1;ram[19][39]=1;ram[19][40]=0;ram[19][41]=1;ram[19][42]=0;ram[19][43]=1;ram[19][44]=0;ram[19][45]=1;ram[19][46]=1;ram[19][47]=1;ram[19][48]=1;ram[19][49]=0;ram[19][50]=1;ram[19][51]=1;ram[19][52]=0;ram[19][53]=0;ram[19][54]=0;ram[19][55]=0;ram[19][56]=1;ram[19][57]=0;ram[19][58]=1;ram[19][59]=1;ram[19][60]=0;ram[19][61]=0;ram[19][62]=1;ram[19][63]=0;ram[19][64]=0;ram[19][65]=0;ram[19][66]=1;ram[19][67]=1;ram[19][68]=1;ram[19][69]=1;ram[19][70]=1;ram[19][71]=1;ram[19][72]=1;ram[19][73]=1;ram[19][74]=1;ram[19][75]=1;ram[19][76]=1;ram[19][77]=0;ram[19][78]=1;ram[19][79]=1;ram[19][80]=1;ram[19][81]=1;ram[19][82]=1;ram[19][83]=1;ram[19][84]=1;ram[19][85]=1;ram[19][86]=0;ram[19][87]=1;ram[19][88]=1;ram[19][89]=1;ram[19][90]=1;ram[19][91]=1;ram[19][92]=1;ram[19][93]=1;ram[19][94]=1;ram[19][95]=0;ram[19][96]=1;ram[19][97]=1;ram[19][98]=0;ram[19][99]=1;ram[19][100]=1;ram[19][101]=1;ram[19][102]=1;ram[19][103]=0;ram[19][104]=1;ram[19][105]=1;ram[19][106]=1;ram[19][107]=0;ram[19][108]=1;ram[19][109]=0;ram[19][110]=0;ram[19][111]=1;ram[19][112]=1;ram[19][113]=1;ram[19][114]=1;ram[19][115]=1;ram[19][116]=0;ram[19][117]=0;ram[19][118]=1;ram[19][119]=1;ram[19][120]=0;ram[19][121]=0;ram[19][122]=1;ram[19][123]=1;ram[19][124]=1;ram[19][125]=1;ram[19][126]=1;ram[19][127]=0;ram[19][128]=1;ram[19][129]=0;ram[19][130]=1;ram[19][131]=1;ram[19][132]=0;ram[19][133]=0;ram[19][134]=1;ram[19][135]=1;ram[19][136]=0;
        ram[20][0]=1;ram[20][1]=1;ram[20][2]=1;ram[20][3]=1;ram[20][4]=1;ram[20][5]=1;ram[20][6]=1;ram[20][7]=1;ram[20][8]=0;ram[20][9]=1;ram[20][10]=1;ram[20][11]=1;ram[20][12]=1;ram[20][13]=1;ram[20][14]=0;ram[20][15]=1;ram[20][16]=1;ram[20][17]=1;ram[20][18]=1;ram[20][19]=0;ram[20][20]=1;ram[20][21]=0;ram[20][22]=0;ram[20][23]=1;ram[20][24]=1;ram[20][25]=1;ram[20][26]=1;ram[20][27]=1;ram[20][28]=0;ram[20][29]=0;ram[20][30]=1;ram[20][31]=0;ram[20][32]=1;ram[20][33]=1;ram[20][34]=1;ram[20][35]=1;ram[20][36]=1;ram[20][37]=1;ram[20][38]=0;ram[20][39]=1;ram[20][40]=1;ram[20][41]=1;ram[20][42]=0;ram[20][43]=0;ram[20][44]=1;ram[20][45]=1;ram[20][46]=0;ram[20][47]=1;ram[20][48]=0;ram[20][49]=1;ram[20][50]=0;ram[20][51]=1;ram[20][52]=0;ram[20][53]=1;ram[20][54]=1;ram[20][55]=0;ram[20][56]=0;ram[20][57]=1;ram[20][58]=1;ram[20][59]=1;ram[20][60]=0;ram[20][61]=1;ram[20][62]=1;ram[20][63]=1;ram[20][64]=0;ram[20][65]=1;ram[20][66]=1;ram[20][67]=1;ram[20][68]=1;ram[20][69]=0;ram[20][70]=1;ram[20][71]=0;ram[20][72]=1;ram[20][73]=1;ram[20][74]=0;ram[20][75]=1;ram[20][76]=1;ram[20][77]=1;ram[20][78]=0;ram[20][79]=0;ram[20][80]=0;ram[20][81]=1;ram[20][82]=1;ram[20][83]=0;ram[20][84]=0;ram[20][85]=1;ram[20][86]=0;ram[20][87]=1;ram[20][88]=1;ram[20][89]=1;ram[20][90]=0;ram[20][91]=0;ram[20][92]=0;ram[20][93]=1;ram[20][94]=0;ram[20][95]=1;ram[20][96]=1;ram[20][97]=1;ram[20][98]=1;ram[20][99]=1;ram[20][100]=1;ram[20][101]=0;ram[20][102]=1;ram[20][103]=1;ram[20][104]=0;ram[20][105]=0;ram[20][106]=1;ram[20][107]=0;ram[20][108]=1;ram[20][109]=0;ram[20][110]=1;ram[20][111]=1;ram[20][112]=1;ram[20][113]=0;ram[20][114]=0;ram[20][115]=1;ram[20][116]=1;ram[20][117]=0;ram[20][118]=1;ram[20][119]=1;ram[20][120]=1;ram[20][121]=1;ram[20][122]=0;ram[20][123]=1;ram[20][124]=0;ram[20][125]=1;ram[20][126]=0;ram[20][127]=1;ram[20][128]=1;ram[20][129]=0;ram[20][130]=0;ram[20][131]=0;ram[20][132]=1;ram[20][133]=1;ram[20][134]=1;ram[20][135]=0;ram[20][136]=1;
        ram[21][0]=1;ram[21][1]=1;ram[21][2]=1;ram[21][3]=0;ram[21][4]=1;ram[21][5]=1;ram[21][6]=1;ram[21][7]=1;ram[21][8]=0;ram[21][9]=1;ram[21][10]=0;ram[21][11]=1;ram[21][12]=0;ram[21][13]=1;ram[21][14]=0;ram[21][15]=1;ram[21][16]=1;ram[21][17]=1;ram[21][18]=1;ram[21][19]=0;ram[21][20]=0;ram[21][21]=0;ram[21][22]=1;ram[21][23]=0;ram[21][24]=1;ram[21][25]=1;ram[21][26]=0;ram[21][27]=1;ram[21][28]=1;ram[21][29]=0;ram[21][30]=0;ram[21][31]=0;ram[21][32]=0;ram[21][33]=0;ram[21][34]=1;ram[21][35]=1;ram[21][36]=0;ram[21][37]=0;ram[21][38]=1;ram[21][39]=0;ram[21][40]=0;ram[21][41]=0;ram[21][42]=0;ram[21][43]=1;ram[21][44]=1;ram[21][45]=1;ram[21][46]=1;ram[21][47]=1;ram[21][48]=0;ram[21][49]=1;ram[21][50]=1;ram[21][51]=0;ram[21][52]=0;ram[21][53]=1;ram[21][54]=1;ram[21][55]=1;ram[21][56]=1;ram[21][57]=1;ram[21][58]=0;ram[21][59]=0;ram[21][60]=1;ram[21][61]=0;ram[21][62]=0;ram[21][63]=1;ram[21][64]=0;ram[21][65]=0;ram[21][66]=1;ram[21][67]=0;ram[21][68]=1;ram[21][69]=1;ram[21][70]=1;ram[21][71]=0;ram[21][72]=1;ram[21][73]=1;ram[21][74]=0;ram[21][75]=1;ram[21][76]=0;ram[21][77]=1;ram[21][78]=1;ram[21][79]=1;ram[21][80]=1;ram[21][81]=1;ram[21][82]=1;ram[21][83]=1;ram[21][84]=0;ram[21][85]=0;ram[21][86]=0;ram[21][87]=1;ram[21][88]=1;ram[21][89]=0;ram[21][90]=1;ram[21][91]=1;ram[21][92]=1;ram[21][93]=1;ram[21][94]=0;ram[21][95]=1;ram[21][96]=1;ram[21][97]=1;ram[21][98]=0;ram[21][99]=1;ram[21][100]=1;ram[21][101]=0;ram[21][102]=0;ram[21][103]=1;ram[21][104]=1;ram[21][105]=0;ram[21][106]=1;ram[21][107]=1;ram[21][108]=1;ram[21][109]=1;ram[21][110]=0;ram[21][111]=0;ram[21][112]=1;ram[21][113]=0;ram[21][114]=1;ram[21][115]=1;ram[21][116]=1;ram[21][117]=0;ram[21][118]=1;ram[21][119]=1;ram[21][120]=1;ram[21][121]=1;ram[21][122]=1;ram[21][123]=1;ram[21][124]=1;ram[21][125]=1;ram[21][126]=1;ram[21][127]=1;ram[21][128]=1;ram[21][129]=1;ram[21][130]=1;ram[21][131]=1;ram[21][132]=0;ram[21][133]=1;ram[21][134]=1;ram[21][135]=0;ram[21][136]=1;
        ram[22][0]=1;ram[22][1]=1;ram[22][2]=1;ram[22][3]=1;ram[22][4]=1;ram[22][5]=1;ram[22][6]=1;ram[22][7]=1;ram[22][8]=1;ram[22][9]=0;ram[22][10]=1;ram[22][11]=1;ram[22][12]=1;ram[22][13]=1;ram[22][14]=0;ram[22][15]=1;ram[22][16]=1;ram[22][17]=0;ram[22][18]=1;ram[22][19]=0;ram[22][20]=1;ram[22][21]=1;ram[22][22]=1;ram[22][23]=1;ram[22][24]=1;ram[22][25]=1;ram[22][26]=0;ram[22][27]=1;ram[22][28]=1;ram[22][29]=0;ram[22][30]=0;ram[22][31]=1;ram[22][32]=1;ram[22][33]=1;ram[22][34]=0;ram[22][35]=1;ram[22][36]=1;ram[22][37]=0;ram[22][38]=1;ram[22][39]=0;ram[22][40]=1;ram[22][41]=1;ram[22][42]=1;ram[22][43]=1;ram[22][44]=1;ram[22][45]=0;ram[22][46]=1;ram[22][47]=0;ram[22][48]=1;ram[22][49]=0;ram[22][50]=0;ram[22][51]=1;ram[22][52]=1;ram[22][53]=1;ram[22][54]=1;ram[22][55]=1;ram[22][56]=0;ram[22][57]=0;ram[22][58]=1;ram[22][59]=1;ram[22][60]=1;ram[22][61]=0;ram[22][62]=1;ram[22][63]=1;ram[22][64]=1;ram[22][65]=1;ram[22][66]=0;ram[22][67]=1;ram[22][68]=1;ram[22][69]=1;ram[22][70]=1;ram[22][71]=1;ram[22][72]=1;ram[22][73]=1;ram[22][74]=1;ram[22][75]=1;ram[22][76]=0;ram[22][77]=1;ram[22][78]=0;ram[22][79]=0;ram[22][80]=0;ram[22][81]=1;ram[22][82]=1;ram[22][83]=1;ram[22][84]=1;ram[22][85]=0;ram[22][86]=0;ram[22][87]=1;ram[22][88]=1;ram[22][89]=1;ram[22][90]=1;ram[22][91]=0;ram[22][92]=0;ram[22][93]=0;ram[22][94]=1;ram[22][95]=0;ram[22][96]=1;ram[22][97]=0;ram[22][98]=0;ram[22][99]=1;ram[22][100]=0;ram[22][101]=0;ram[22][102]=0;ram[22][103]=0;ram[22][104]=1;ram[22][105]=0;ram[22][106]=0;ram[22][107]=1;ram[22][108]=0;ram[22][109]=0;ram[22][110]=1;ram[22][111]=0;ram[22][112]=0;ram[22][113]=1;ram[22][114]=1;ram[22][115]=0;ram[22][116]=1;ram[22][117]=1;ram[22][118]=1;ram[22][119]=1;ram[22][120]=1;ram[22][121]=1;ram[22][122]=1;ram[22][123]=1;ram[22][124]=0;ram[22][125]=1;ram[22][126]=1;ram[22][127]=1;ram[22][128]=1;ram[22][129]=0;ram[22][130]=0;ram[22][131]=1;ram[22][132]=1;ram[22][133]=0;ram[22][134]=1;ram[22][135]=1;ram[22][136]=0;
        ram[23][0]=1;ram[23][1]=1;ram[23][2]=0;ram[23][3]=1;ram[23][4]=0;ram[23][5]=1;ram[23][6]=0;ram[23][7]=0;ram[23][8]=1;ram[23][9]=0;ram[23][10]=1;ram[23][11]=1;ram[23][12]=1;ram[23][13]=1;ram[23][14]=1;ram[23][15]=0;ram[23][16]=0;ram[23][17]=1;ram[23][18]=1;ram[23][19]=1;ram[23][20]=1;ram[23][21]=0;ram[23][22]=0;ram[23][23]=1;ram[23][24]=0;ram[23][25]=0;ram[23][26]=1;ram[23][27]=1;ram[23][28]=1;ram[23][29]=1;ram[23][30]=1;ram[23][31]=0;ram[23][32]=1;ram[23][33]=0;ram[23][34]=1;ram[23][35]=0;ram[23][36]=1;ram[23][37]=0;ram[23][38]=1;ram[23][39]=1;ram[23][40]=0;ram[23][41]=1;ram[23][42]=0;ram[23][43]=1;ram[23][44]=0;ram[23][45]=0;ram[23][46]=1;ram[23][47]=1;ram[23][48]=0;ram[23][49]=1;ram[23][50]=1;ram[23][51]=0;ram[23][52]=1;ram[23][53]=0;ram[23][54]=1;ram[23][55]=0;ram[23][56]=1;ram[23][57]=0;ram[23][58]=0;ram[23][59]=1;ram[23][60]=0;ram[23][61]=0;ram[23][62]=0;ram[23][63]=0;ram[23][64]=1;ram[23][65]=0;ram[23][66]=0;ram[23][67]=1;ram[23][68]=1;ram[23][69]=1;ram[23][70]=1;ram[23][71]=1;ram[23][72]=1;ram[23][73]=1;ram[23][74]=0;ram[23][75]=1;ram[23][76]=1;ram[23][77]=0;ram[23][78]=1;ram[23][79]=0;ram[23][80]=1;ram[23][81]=1;ram[23][82]=1;ram[23][83]=1;ram[23][84]=1;ram[23][85]=1;ram[23][86]=1;ram[23][87]=1;ram[23][88]=1;ram[23][89]=1;ram[23][90]=1;ram[23][91]=1;ram[23][92]=0;ram[23][93]=0;ram[23][94]=1;ram[23][95]=1;ram[23][96]=1;ram[23][97]=0;ram[23][98]=1;ram[23][99]=0;ram[23][100]=1;ram[23][101]=0;ram[23][102]=1;ram[23][103]=0;ram[23][104]=1;ram[23][105]=0;ram[23][106]=0;ram[23][107]=1;ram[23][108]=0;ram[23][109]=0;ram[23][110]=0;ram[23][111]=1;ram[23][112]=0;ram[23][113]=0;ram[23][114]=0;ram[23][115]=1;ram[23][116]=1;ram[23][117]=1;ram[23][118]=1;ram[23][119]=1;ram[23][120]=0;ram[23][121]=1;ram[23][122]=1;ram[23][123]=0;ram[23][124]=0;ram[23][125]=1;ram[23][126]=1;ram[23][127]=1;ram[23][128]=0;ram[23][129]=1;ram[23][130]=0;ram[23][131]=0;ram[23][132]=1;ram[23][133]=0;ram[23][134]=1;ram[23][135]=1;ram[23][136]=0;
        ram[24][0]=0;ram[24][1]=0;ram[24][2]=1;ram[24][3]=1;ram[24][4]=0;ram[24][5]=1;ram[24][6]=1;ram[24][7]=0;ram[24][8]=1;ram[24][9]=0;ram[24][10]=0;ram[24][11]=1;ram[24][12]=1;ram[24][13]=1;ram[24][14]=1;ram[24][15]=0;ram[24][16]=1;ram[24][17]=1;ram[24][18]=1;ram[24][19]=1;ram[24][20]=1;ram[24][21]=0;ram[24][22]=0;ram[24][23]=1;ram[24][24]=1;ram[24][25]=0;ram[24][26]=1;ram[24][27]=1;ram[24][28]=1;ram[24][29]=1;ram[24][30]=0;ram[24][31]=1;ram[24][32]=0;ram[24][33]=1;ram[24][34]=1;ram[24][35]=0;ram[24][36]=1;ram[24][37]=1;ram[24][38]=1;ram[24][39]=1;ram[24][40]=0;ram[24][41]=1;ram[24][42]=1;ram[24][43]=0;ram[24][44]=1;ram[24][45]=0;ram[24][46]=1;ram[24][47]=1;ram[24][48]=0;ram[24][49]=1;ram[24][50]=1;ram[24][51]=0;ram[24][52]=0;ram[24][53]=1;ram[24][54]=1;ram[24][55]=1;ram[24][56]=1;ram[24][57]=0;ram[24][58]=1;ram[24][59]=1;ram[24][60]=1;ram[24][61]=1;ram[24][62]=0;ram[24][63]=1;ram[24][64]=1;ram[24][65]=1;ram[24][66]=0;ram[24][67]=1;ram[24][68]=0;ram[24][69]=1;ram[24][70]=1;ram[24][71]=1;ram[24][72]=1;ram[24][73]=0;ram[24][74]=1;ram[24][75]=1;ram[24][76]=1;ram[24][77]=0;ram[24][78]=1;ram[24][79]=0;ram[24][80]=0;ram[24][81]=0;ram[24][82]=1;ram[24][83]=0;ram[24][84]=0;ram[24][85]=0;ram[24][86]=0;ram[24][87]=0;ram[24][88]=1;ram[24][89]=1;ram[24][90]=0;ram[24][91]=1;ram[24][92]=0;ram[24][93]=1;ram[24][94]=1;ram[24][95]=0;ram[24][96]=0;ram[24][97]=1;ram[24][98]=0;ram[24][99]=1;ram[24][100]=0;ram[24][101]=1;ram[24][102]=1;ram[24][103]=0;ram[24][104]=0;ram[24][105]=1;ram[24][106]=1;ram[24][107]=1;ram[24][108]=0;ram[24][109]=0;ram[24][110]=1;ram[24][111]=1;ram[24][112]=1;ram[24][113]=1;ram[24][114]=1;ram[24][115]=1;ram[24][116]=0;ram[24][117]=0;ram[24][118]=1;ram[24][119]=0;ram[24][120]=1;ram[24][121]=1;ram[24][122]=1;ram[24][123]=1;ram[24][124]=1;ram[24][125]=1;ram[24][126]=0;ram[24][127]=0;ram[24][128]=0;ram[24][129]=0;ram[24][130]=1;ram[24][131]=0;ram[24][132]=0;ram[24][133]=1;ram[24][134]=1;ram[24][135]=1;ram[24][136]=0;
        ram[25][0]=1;ram[25][1]=1;ram[25][2]=1;ram[25][3]=0;ram[25][4]=0;ram[25][5]=1;ram[25][6]=1;ram[25][7]=1;ram[25][8]=1;ram[25][9]=1;ram[25][10]=0;ram[25][11]=1;ram[25][12]=0;ram[25][13]=1;ram[25][14]=1;ram[25][15]=1;ram[25][16]=0;ram[25][17]=0;ram[25][18]=1;ram[25][19]=0;ram[25][20]=0;ram[25][21]=1;ram[25][22]=1;ram[25][23]=1;ram[25][24]=1;ram[25][25]=0;ram[25][26]=1;ram[25][27]=0;ram[25][28]=1;ram[25][29]=0;ram[25][30]=1;ram[25][31]=1;ram[25][32]=1;ram[25][33]=0;ram[25][34]=1;ram[25][35]=1;ram[25][36]=0;ram[25][37]=1;ram[25][38]=0;ram[25][39]=0;ram[25][40]=0;ram[25][41]=1;ram[25][42]=0;ram[25][43]=0;ram[25][44]=0;ram[25][45]=0;ram[25][46]=1;ram[25][47]=1;ram[25][48]=1;ram[25][49]=1;ram[25][50]=1;ram[25][51]=0;ram[25][52]=1;ram[25][53]=1;ram[25][54]=0;ram[25][55]=0;ram[25][56]=1;ram[25][57]=1;ram[25][58]=1;ram[25][59]=0;ram[25][60]=1;ram[25][61]=1;ram[25][62]=0;ram[25][63]=1;ram[25][64]=1;ram[25][65]=1;ram[25][66]=0;ram[25][67]=1;ram[25][68]=1;ram[25][69]=1;ram[25][70]=0;ram[25][71]=1;ram[25][72]=1;ram[25][73]=0;ram[25][74]=0;ram[25][75]=1;ram[25][76]=0;ram[25][77]=0;ram[25][78]=0;ram[25][79]=1;ram[25][80]=1;ram[25][81]=0;ram[25][82]=0;ram[25][83]=0;ram[25][84]=0;ram[25][85]=1;ram[25][86]=0;ram[25][87]=1;ram[25][88]=1;ram[25][89]=1;ram[25][90]=1;ram[25][91]=1;ram[25][92]=1;ram[25][93]=1;ram[25][94]=0;ram[25][95]=1;ram[25][96]=1;ram[25][97]=0;ram[25][98]=0;ram[25][99]=0;ram[25][100]=1;ram[25][101]=0;ram[25][102]=0;ram[25][103]=1;ram[25][104]=0;ram[25][105]=1;ram[25][106]=0;ram[25][107]=1;ram[25][108]=1;ram[25][109]=0;ram[25][110]=0;ram[25][111]=1;ram[25][112]=1;ram[25][113]=0;ram[25][114]=0;ram[25][115]=1;ram[25][116]=1;ram[25][117]=0;ram[25][118]=1;ram[25][119]=0;ram[25][120]=0;ram[25][121]=1;ram[25][122]=1;ram[25][123]=1;ram[25][124]=1;ram[25][125]=0;ram[25][126]=1;ram[25][127]=1;ram[25][128]=1;ram[25][129]=1;ram[25][130]=0;ram[25][131]=1;ram[25][132]=1;ram[25][133]=1;ram[25][134]=1;ram[25][135]=1;ram[25][136]=0;
        ram[26][0]=0;ram[26][1]=1;ram[26][2]=0;ram[26][3]=1;ram[26][4]=1;ram[26][5]=0;ram[26][6]=1;ram[26][7]=1;ram[26][8]=1;ram[26][9]=1;ram[26][10]=0;ram[26][11]=1;ram[26][12]=0;ram[26][13]=0;ram[26][14]=1;ram[26][15]=1;ram[26][16]=1;ram[26][17]=1;ram[26][18]=0;ram[26][19]=1;ram[26][20]=1;ram[26][21]=1;ram[26][22]=1;ram[26][23]=1;ram[26][24]=1;ram[26][25]=1;ram[26][26]=0;ram[26][27]=1;ram[26][28]=1;ram[26][29]=1;ram[26][30]=1;ram[26][31]=1;ram[26][32]=1;ram[26][33]=0;ram[26][34]=1;ram[26][35]=0;ram[26][36]=1;ram[26][37]=1;ram[26][38]=1;ram[26][39]=1;ram[26][40]=1;ram[26][41]=1;ram[26][42]=1;ram[26][43]=0;ram[26][44]=1;ram[26][45]=1;ram[26][46]=1;ram[26][47]=0;ram[26][48]=1;ram[26][49]=1;ram[26][50]=1;ram[26][51]=1;ram[26][52]=1;ram[26][53]=0;ram[26][54]=1;ram[26][55]=1;ram[26][56]=1;ram[26][57]=0;ram[26][58]=1;ram[26][59]=0;ram[26][60]=1;ram[26][61]=0;ram[26][62]=0;ram[26][63]=0;ram[26][64]=0;ram[26][65]=0;ram[26][66]=1;ram[26][67]=1;ram[26][68]=1;ram[26][69]=1;ram[26][70]=0;ram[26][71]=0;ram[26][72]=0;ram[26][73]=0;ram[26][74]=1;ram[26][75]=0;ram[26][76]=0;ram[26][77]=1;ram[26][78]=0;ram[26][79]=1;ram[26][80]=1;ram[26][81]=1;ram[26][82]=0;ram[26][83]=1;ram[26][84]=1;ram[26][85]=1;ram[26][86]=1;ram[26][87]=1;ram[26][88]=1;ram[26][89]=0;ram[26][90]=0;ram[26][91]=0;ram[26][92]=1;ram[26][93]=1;ram[26][94]=1;ram[26][95]=0;ram[26][96]=0;ram[26][97]=1;ram[26][98]=1;ram[26][99]=0;ram[26][100]=1;ram[26][101]=1;ram[26][102]=0;ram[26][103]=1;ram[26][104]=1;ram[26][105]=1;ram[26][106]=0;ram[26][107]=0;ram[26][108]=0;ram[26][109]=1;ram[26][110]=1;ram[26][111]=1;ram[26][112]=1;ram[26][113]=1;ram[26][114]=1;ram[26][115]=1;ram[26][116]=1;ram[26][117]=0;ram[26][118]=1;ram[26][119]=1;ram[26][120]=1;ram[26][121]=1;ram[26][122]=1;ram[26][123]=1;ram[26][124]=0;ram[26][125]=0;ram[26][126]=0;ram[26][127]=1;ram[26][128]=1;ram[26][129]=1;ram[26][130]=0;ram[26][131]=1;ram[26][132]=1;ram[26][133]=1;ram[26][134]=1;ram[26][135]=0;ram[26][136]=0;
        ram[27][0]=1;ram[27][1]=0;ram[27][2]=0;ram[27][3]=1;ram[27][4]=1;ram[27][5]=1;ram[27][6]=0;ram[27][7]=1;ram[27][8]=1;ram[27][9]=1;ram[27][10]=0;ram[27][11]=1;ram[27][12]=0;ram[27][13]=0;ram[27][14]=0;ram[27][15]=1;ram[27][16]=1;ram[27][17]=0;ram[27][18]=0;ram[27][19]=1;ram[27][20]=0;ram[27][21]=1;ram[27][22]=0;ram[27][23]=1;ram[27][24]=1;ram[27][25]=0;ram[27][26]=1;ram[27][27]=1;ram[27][28]=1;ram[27][29]=0;ram[27][30]=1;ram[27][31]=0;ram[27][32]=0;ram[27][33]=0;ram[27][34]=0;ram[27][35]=1;ram[27][36]=0;ram[27][37]=0;ram[27][38]=0;ram[27][39]=1;ram[27][40]=0;ram[27][41]=1;ram[27][42]=1;ram[27][43]=0;ram[27][44]=1;ram[27][45]=1;ram[27][46]=1;ram[27][47]=1;ram[27][48]=0;ram[27][49]=1;ram[27][50]=1;ram[27][51]=0;ram[27][52]=1;ram[27][53]=0;ram[27][54]=0;ram[27][55]=1;ram[27][56]=0;ram[27][57]=1;ram[27][58]=1;ram[27][59]=1;ram[27][60]=0;ram[27][61]=1;ram[27][62]=0;ram[27][63]=0;ram[27][64]=1;ram[27][65]=1;ram[27][66]=1;ram[27][67]=1;ram[27][68]=0;ram[27][69]=1;ram[27][70]=1;ram[27][71]=0;ram[27][72]=1;ram[27][73]=0;ram[27][74]=1;ram[27][75]=1;ram[27][76]=1;ram[27][77]=1;ram[27][78]=1;ram[27][79]=1;ram[27][80]=1;ram[27][81]=0;ram[27][82]=0;ram[27][83]=1;ram[27][84]=1;ram[27][85]=1;ram[27][86]=1;ram[27][87]=1;ram[27][88]=1;ram[27][89]=1;ram[27][90]=1;ram[27][91]=1;ram[27][92]=1;ram[27][93]=1;ram[27][94]=0;ram[27][95]=0;ram[27][96]=0;ram[27][97]=1;ram[27][98]=1;ram[27][99]=1;ram[27][100]=0;ram[27][101]=1;ram[27][102]=0;ram[27][103]=1;ram[27][104]=1;ram[27][105]=1;ram[27][106]=0;ram[27][107]=1;ram[27][108]=1;ram[27][109]=0;ram[27][110]=0;ram[27][111]=0;ram[27][112]=1;ram[27][113]=1;ram[27][114]=1;ram[27][115]=1;ram[27][116]=1;ram[27][117]=1;ram[27][118]=1;ram[27][119]=0;ram[27][120]=0;ram[27][121]=1;ram[27][122]=1;ram[27][123]=1;ram[27][124]=0;ram[27][125]=1;ram[27][126]=1;ram[27][127]=1;ram[27][128]=1;ram[27][129]=0;ram[27][130]=0;ram[27][131]=1;ram[27][132]=1;ram[27][133]=0;ram[27][134]=0;ram[27][135]=1;ram[27][136]=1;
        ram[28][0]=1;ram[28][1]=0;ram[28][2]=0;ram[28][3]=1;ram[28][4]=0;ram[28][5]=1;ram[28][6]=1;ram[28][7]=1;ram[28][8]=1;ram[28][9]=0;ram[28][10]=1;ram[28][11]=1;ram[28][12]=1;ram[28][13]=1;ram[28][14]=0;ram[28][15]=0;ram[28][16]=1;ram[28][17]=0;ram[28][18]=0;ram[28][19]=1;ram[28][20]=1;ram[28][21]=0;ram[28][22]=0;ram[28][23]=1;ram[28][24]=0;ram[28][25]=1;ram[28][26]=1;ram[28][27]=0;ram[28][28]=1;ram[28][29]=1;ram[28][30]=1;ram[28][31]=1;ram[28][32]=1;ram[28][33]=0;ram[28][34]=1;ram[28][35]=1;ram[28][36]=0;ram[28][37]=1;ram[28][38]=0;ram[28][39]=0;ram[28][40]=1;ram[28][41]=0;ram[28][42]=0;ram[28][43]=1;ram[28][44]=1;ram[28][45]=0;ram[28][46]=1;ram[28][47]=1;ram[28][48]=1;ram[28][49]=0;ram[28][50]=0;ram[28][51]=0;ram[28][52]=1;ram[28][53]=1;ram[28][54]=1;ram[28][55]=1;ram[28][56]=1;ram[28][57]=1;ram[28][58]=1;ram[28][59]=0;ram[28][60]=1;ram[28][61]=1;ram[28][62]=0;ram[28][63]=0;ram[28][64]=0;ram[28][65]=0;ram[28][66]=1;ram[28][67]=1;ram[28][68]=1;ram[28][69]=1;ram[28][70]=1;ram[28][71]=1;ram[28][72]=0;ram[28][73]=1;ram[28][74]=1;ram[28][75]=1;ram[28][76]=0;ram[28][77]=1;ram[28][78]=1;ram[28][79]=0;ram[28][80]=1;ram[28][81]=1;ram[28][82]=0;ram[28][83]=1;ram[28][84]=1;ram[28][85]=1;ram[28][86]=1;ram[28][87]=1;ram[28][88]=1;ram[28][89]=1;ram[28][90]=1;ram[28][91]=1;ram[28][92]=1;ram[28][93]=0;ram[28][94]=0;ram[28][95]=1;ram[28][96]=1;ram[28][97]=0;ram[28][98]=1;ram[28][99]=1;ram[28][100]=1;ram[28][101]=0;ram[28][102]=1;ram[28][103]=1;ram[28][104]=1;ram[28][105]=1;ram[28][106]=0;ram[28][107]=1;ram[28][108]=1;ram[28][109]=0;ram[28][110]=1;ram[28][111]=0;ram[28][112]=1;ram[28][113]=0;ram[28][114]=0;ram[28][115]=0;ram[28][116]=1;ram[28][117]=1;ram[28][118]=0;ram[28][119]=1;ram[28][120]=1;ram[28][121]=0;ram[28][122]=1;ram[28][123]=1;ram[28][124]=1;ram[28][125]=0;ram[28][126]=0;ram[28][127]=0;ram[28][128]=1;ram[28][129]=1;ram[28][130]=1;ram[28][131]=1;ram[28][132]=1;ram[28][133]=1;ram[28][134]=0;ram[28][135]=0;ram[28][136]=1;
        ram[29][0]=1;ram[29][1]=0;ram[29][2]=1;ram[29][3]=1;ram[29][4]=1;ram[29][5]=1;ram[29][6]=0;ram[29][7]=0;ram[29][8]=0;ram[29][9]=1;ram[29][10]=1;ram[29][11]=1;ram[29][12]=0;ram[29][13]=0;ram[29][14]=0;ram[29][15]=0;ram[29][16]=1;ram[29][17]=1;ram[29][18]=0;ram[29][19]=1;ram[29][20]=1;ram[29][21]=1;ram[29][22]=0;ram[29][23]=0;ram[29][24]=0;ram[29][25]=1;ram[29][26]=1;ram[29][27]=1;ram[29][28]=1;ram[29][29]=1;ram[29][30]=1;ram[29][31]=0;ram[29][32]=1;ram[29][33]=1;ram[29][34]=1;ram[29][35]=0;ram[29][36]=1;ram[29][37]=0;ram[29][38]=1;ram[29][39]=0;ram[29][40]=1;ram[29][41]=1;ram[29][42]=0;ram[29][43]=1;ram[29][44]=1;ram[29][45]=1;ram[29][46]=1;ram[29][47]=1;ram[29][48]=1;ram[29][49]=0;ram[29][50]=1;ram[29][51]=1;ram[29][52]=1;ram[29][53]=1;ram[29][54]=1;ram[29][55]=1;ram[29][56]=0;ram[29][57]=0;ram[29][58]=1;ram[29][59]=0;ram[29][60]=0;ram[29][61]=0;ram[29][62]=0;ram[29][63]=1;ram[29][64]=1;ram[29][65]=1;ram[29][66]=1;ram[29][67]=0;ram[29][68]=1;ram[29][69]=0;ram[29][70]=0;ram[29][71]=1;ram[29][72]=0;ram[29][73]=0;ram[29][74]=1;ram[29][75]=0;ram[29][76]=0;ram[29][77]=0;ram[29][78]=1;ram[29][79]=1;ram[29][80]=0;ram[29][81]=1;ram[29][82]=1;ram[29][83]=1;ram[29][84]=1;ram[29][85]=1;ram[29][86]=1;ram[29][87]=1;ram[29][88]=0;ram[29][89]=0;ram[29][90]=1;ram[29][91]=0;ram[29][92]=1;ram[29][93]=1;ram[29][94]=1;ram[29][95]=0;ram[29][96]=1;ram[29][97]=1;ram[29][98]=1;ram[29][99]=1;ram[29][100]=1;ram[29][101]=1;ram[29][102]=1;ram[29][103]=1;ram[29][104]=1;ram[29][105]=1;ram[29][106]=1;ram[29][107]=1;ram[29][108]=1;ram[29][109]=0;ram[29][110]=1;ram[29][111]=1;ram[29][112]=1;ram[29][113]=1;ram[29][114]=1;ram[29][115]=1;ram[29][116]=1;ram[29][117]=1;ram[29][118]=1;ram[29][119]=1;ram[29][120]=0;ram[29][121]=1;ram[29][122]=1;ram[29][123]=0;ram[29][124]=1;ram[29][125]=1;ram[29][126]=1;ram[29][127]=1;ram[29][128]=1;ram[29][129]=1;ram[29][130]=0;ram[29][131]=0;ram[29][132]=0;ram[29][133]=1;ram[29][134]=1;ram[29][135]=0;ram[29][136]=1;
        ram[30][0]=0;ram[30][1]=1;ram[30][2]=0;ram[30][3]=0;ram[30][4]=1;ram[30][5]=1;ram[30][6]=1;ram[30][7]=1;ram[30][8]=0;ram[30][9]=1;ram[30][10]=0;ram[30][11]=0;ram[30][12]=0;ram[30][13]=1;ram[30][14]=0;ram[30][15]=1;ram[30][16]=1;ram[30][17]=0;ram[30][18]=1;ram[30][19]=1;ram[30][20]=1;ram[30][21]=1;ram[30][22]=1;ram[30][23]=1;ram[30][24]=0;ram[30][25]=1;ram[30][26]=1;ram[30][27]=1;ram[30][28]=1;ram[30][29]=1;ram[30][30]=1;ram[30][31]=0;ram[30][32]=1;ram[30][33]=1;ram[30][34]=1;ram[30][35]=0;ram[30][36]=1;ram[30][37]=1;ram[30][38]=1;ram[30][39]=1;ram[30][40]=1;ram[30][41]=1;ram[30][42]=0;ram[30][43]=0;ram[30][44]=1;ram[30][45]=0;ram[30][46]=1;ram[30][47]=1;ram[30][48]=1;ram[30][49]=1;ram[30][50]=1;ram[30][51]=1;ram[30][52]=1;ram[30][53]=1;ram[30][54]=0;ram[30][55]=1;ram[30][56]=0;ram[30][57]=1;ram[30][58]=1;ram[30][59]=1;ram[30][60]=1;ram[30][61]=1;ram[30][62]=0;ram[30][63]=0;ram[30][64]=1;ram[30][65]=0;ram[30][66]=1;ram[30][67]=0;ram[30][68]=0;ram[30][69]=1;ram[30][70]=0;ram[30][71]=0;ram[30][72]=1;ram[30][73]=1;ram[30][74]=0;ram[30][75]=1;ram[30][76]=1;ram[30][77]=1;ram[30][78]=1;ram[30][79]=1;ram[30][80]=0;ram[30][81]=1;ram[30][82]=0;ram[30][83]=0;ram[30][84]=1;ram[30][85]=0;ram[30][86]=0;ram[30][87]=0;ram[30][88]=0;ram[30][89]=1;ram[30][90]=1;ram[30][91]=1;ram[30][92]=1;ram[30][93]=0;ram[30][94]=0;ram[30][95]=0;ram[30][96]=0;ram[30][97]=1;ram[30][98]=1;ram[30][99]=0;ram[30][100]=1;ram[30][101]=1;ram[30][102]=1;ram[30][103]=0;ram[30][104]=1;ram[30][105]=1;ram[30][106]=1;ram[30][107]=1;ram[30][108]=1;ram[30][109]=1;ram[30][110]=1;ram[30][111]=1;ram[30][112]=1;ram[30][113]=1;ram[30][114]=1;ram[30][115]=0;ram[30][116]=1;ram[30][117]=0;ram[30][118]=0;ram[30][119]=0;ram[30][120]=1;ram[30][121]=1;ram[30][122]=1;ram[30][123]=1;ram[30][124]=0;ram[30][125]=1;ram[30][126]=0;ram[30][127]=1;ram[30][128]=1;ram[30][129]=0;ram[30][130]=0;ram[30][131]=1;ram[30][132]=1;ram[30][133]=1;ram[30][134]=1;ram[30][135]=0;ram[30][136]=0;
        ram[31][0]=1;ram[31][1]=0;ram[31][2]=1;ram[31][3]=1;ram[31][4]=1;ram[31][5]=0;ram[31][6]=1;ram[31][7]=0;ram[31][8]=0;ram[31][9]=0;ram[31][10]=0;ram[31][11]=1;ram[31][12]=1;ram[31][13]=1;ram[31][14]=1;ram[31][15]=0;ram[31][16]=0;ram[31][17]=1;ram[31][18]=0;ram[31][19]=1;ram[31][20]=1;ram[31][21]=1;ram[31][22]=0;ram[31][23]=1;ram[31][24]=1;ram[31][25]=1;ram[31][26]=1;ram[31][27]=1;ram[31][28]=1;ram[31][29]=0;ram[31][30]=1;ram[31][31]=0;ram[31][32]=1;ram[31][33]=1;ram[31][34]=1;ram[31][35]=1;ram[31][36]=1;ram[31][37]=1;ram[31][38]=1;ram[31][39]=1;ram[31][40]=1;ram[31][41]=1;ram[31][42]=1;ram[31][43]=1;ram[31][44]=1;ram[31][45]=1;ram[31][46]=1;ram[31][47]=1;ram[31][48]=1;ram[31][49]=1;ram[31][50]=1;ram[31][51]=1;ram[31][52]=0;ram[31][53]=0;ram[31][54]=0;ram[31][55]=1;ram[31][56]=0;ram[31][57]=0;ram[31][58]=1;ram[31][59]=0;ram[31][60]=1;ram[31][61]=1;ram[31][62]=0;ram[31][63]=1;ram[31][64]=1;ram[31][65]=1;ram[31][66]=1;ram[31][67]=1;ram[31][68]=1;ram[31][69]=1;ram[31][70]=0;ram[31][71]=1;ram[31][72]=1;ram[31][73]=1;ram[31][74]=1;ram[31][75]=1;ram[31][76]=0;ram[31][77]=0;ram[31][78]=1;ram[31][79]=1;ram[31][80]=0;ram[31][81]=0;ram[31][82]=1;ram[31][83]=1;ram[31][84]=1;ram[31][85]=1;ram[31][86]=1;ram[31][87]=0;ram[31][88]=0;ram[31][89]=0;ram[31][90]=1;ram[31][91]=1;ram[31][92]=0;ram[31][93]=1;ram[31][94]=1;ram[31][95]=0;ram[31][96]=1;ram[31][97]=1;ram[31][98]=1;ram[31][99]=0;ram[31][100]=1;ram[31][101]=1;ram[31][102]=1;ram[31][103]=0;ram[31][104]=1;ram[31][105]=0;ram[31][106]=1;ram[31][107]=0;ram[31][108]=0;ram[31][109]=0;ram[31][110]=1;ram[31][111]=0;ram[31][112]=0;ram[31][113]=1;ram[31][114]=1;ram[31][115]=1;ram[31][116]=1;ram[31][117]=1;ram[31][118]=0;ram[31][119]=1;ram[31][120]=1;ram[31][121]=1;ram[31][122]=0;ram[31][123]=0;ram[31][124]=1;ram[31][125]=1;ram[31][126]=1;ram[31][127]=0;ram[31][128]=1;ram[31][129]=1;ram[31][130]=1;ram[31][131]=0;ram[31][132]=1;ram[31][133]=1;ram[31][134]=1;ram[31][135]=1;ram[31][136]=0;
        ram[32][0]=1;ram[32][1]=1;ram[32][2]=0;ram[32][3]=0;ram[32][4]=1;ram[32][5]=0;ram[32][6]=1;ram[32][7]=0;ram[32][8]=0;ram[32][9]=0;ram[32][10]=0;ram[32][11]=0;ram[32][12]=0;ram[32][13]=1;ram[32][14]=1;ram[32][15]=1;ram[32][16]=0;ram[32][17]=1;ram[32][18]=1;ram[32][19]=1;ram[32][20]=1;ram[32][21]=0;ram[32][22]=0;ram[32][23]=1;ram[32][24]=1;ram[32][25]=0;ram[32][26]=1;ram[32][27]=1;ram[32][28]=0;ram[32][29]=0;ram[32][30]=1;ram[32][31]=1;ram[32][32]=0;ram[32][33]=1;ram[32][34]=1;ram[32][35]=1;ram[32][36]=0;ram[32][37]=0;ram[32][38]=0;ram[32][39]=1;ram[32][40]=1;ram[32][41]=1;ram[32][42]=1;ram[32][43]=1;ram[32][44]=0;ram[32][45]=1;ram[32][46]=1;ram[32][47]=0;ram[32][48]=0;ram[32][49]=1;ram[32][50]=0;ram[32][51]=0;ram[32][52]=1;ram[32][53]=1;ram[32][54]=0;ram[32][55]=1;ram[32][56]=1;ram[32][57]=1;ram[32][58]=1;ram[32][59]=1;ram[32][60]=1;ram[32][61]=1;ram[32][62]=1;ram[32][63]=1;ram[32][64]=1;ram[32][65]=1;ram[32][66]=0;ram[32][67]=1;ram[32][68]=1;ram[32][69]=1;ram[32][70]=1;ram[32][71]=1;ram[32][72]=1;ram[32][73]=0;ram[32][74]=0;ram[32][75]=1;ram[32][76]=0;ram[32][77]=1;ram[32][78]=1;ram[32][79]=0;ram[32][80]=1;ram[32][81]=1;ram[32][82]=1;ram[32][83]=1;ram[32][84]=1;ram[32][85]=1;ram[32][86]=1;ram[32][87]=1;ram[32][88]=1;ram[32][89]=1;ram[32][90]=0;ram[32][91]=0;ram[32][92]=0;ram[32][93]=0;ram[32][94]=0;ram[32][95]=1;ram[32][96]=1;ram[32][97]=1;ram[32][98]=0;ram[32][99]=1;ram[32][100]=0;ram[32][101]=1;ram[32][102]=1;ram[32][103]=1;ram[32][104]=1;ram[32][105]=1;ram[32][106]=1;ram[32][107]=1;ram[32][108]=1;ram[32][109]=1;ram[32][110]=1;ram[32][111]=1;ram[32][112]=1;ram[32][113]=1;ram[32][114]=0;ram[32][115]=1;ram[32][116]=1;ram[32][117]=1;ram[32][118]=0;ram[32][119]=1;ram[32][120]=1;ram[32][121]=1;ram[32][122]=0;ram[32][123]=1;ram[32][124]=1;ram[32][125]=1;ram[32][126]=1;ram[32][127]=1;ram[32][128]=1;ram[32][129]=0;ram[32][130]=0;ram[32][131]=1;ram[32][132]=1;ram[32][133]=0;ram[32][134]=1;ram[32][135]=0;ram[32][136]=1;
        ram[33][0]=0;ram[33][1]=1;ram[33][2]=0;ram[33][3]=1;ram[33][4]=1;ram[33][5]=1;ram[33][6]=0;ram[33][7]=0;ram[33][8]=1;ram[33][9]=0;ram[33][10]=0;ram[33][11]=0;ram[33][12]=0;ram[33][13]=1;ram[33][14]=1;ram[33][15]=1;ram[33][16]=1;ram[33][17]=0;ram[33][18]=0;ram[33][19]=1;ram[33][20]=1;ram[33][21]=0;ram[33][22]=1;ram[33][23]=1;ram[33][24]=1;ram[33][25]=0;ram[33][26]=1;ram[33][27]=1;ram[33][28]=1;ram[33][29]=1;ram[33][30]=1;ram[33][31]=1;ram[33][32]=1;ram[33][33]=1;ram[33][34]=1;ram[33][35]=1;ram[33][36]=1;ram[33][37]=1;ram[33][38]=0;ram[33][39]=0;ram[33][40]=1;ram[33][41]=1;ram[33][42]=0;ram[33][43]=0;ram[33][44]=1;ram[33][45]=1;ram[33][46]=0;ram[33][47]=1;ram[33][48]=1;ram[33][49]=1;ram[33][50]=1;ram[33][51]=1;ram[33][52]=1;ram[33][53]=0;ram[33][54]=1;ram[33][55]=0;ram[33][56]=1;ram[33][57]=0;ram[33][58]=1;ram[33][59]=1;ram[33][60]=1;ram[33][61]=0;ram[33][62]=0;ram[33][63]=1;ram[33][64]=1;ram[33][65]=1;ram[33][66]=0;ram[33][67]=1;ram[33][68]=1;ram[33][69]=1;ram[33][70]=1;ram[33][71]=1;ram[33][72]=1;ram[33][73]=0;ram[33][74]=1;ram[33][75]=1;ram[33][76]=1;ram[33][77]=1;ram[33][78]=0;ram[33][79]=0;ram[33][80]=0;ram[33][81]=1;ram[33][82]=1;ram[33][83]=1;ram[33][84]=1;ram[33][85]=1;ram[33][86]=0;ram[33][87]=1;ram[33][88]=0;ram[33][89]=1;ram[33][90]=1;ram[33][91]=1;ram[33][92]=1;ram[33][93]=0;ram[33][94]=0;ram[33][95]=1;ram[33][96]=1;ram[33][97]=1;ram[33][98]=1;ram[33][99]=1;ram[33][100]=1;ram[33][101]=0;ram[33][102]=1;ram[33][103]=0;ram[33][104]=0;ram[33][105]=1;ram[33][106]=1;ram[33][107]=1;ram[33][108]=1;ram[33][109]=1;ram[33][110]=0;ram[33][111]=1;ram[33][112]=1;ram[33][113]=1;ram[33][114]=1;ram[33][115]=1;ram[33][116]=0;ram[33][117]=0;ram[33][118]=1;ram[33][119]=1;ram[33][120]=1;ram[33][121]=1;ram[33][122]=1;ram[33][123]=1;ram[33][124]=0;ram[33][125]=1;ram[33][126]=0;ram[33][127]=1;ram[33][128]=1;ram[33][129]=1;ram[33][130]=1;ram[33][131]=1;ram[33][132]=1;ram[33][133]=1;ram[33][134]=1;ram[33][135]=1;ram[33][136]=0;
        ram[34][0]=1;ram[34][1]=0;ram[34][2]=0;ram[34][3]=1;ram[34][4]=1;ram[34][5]=1;ram[34][6]=1;ram[34][7]=0;ram[34][8]=1;ram[34][9]=1;ram[34][10]=1;ram[34][11]=1;ram[34][12]=0;ram[34][13]=1;ram[34][14]=0;ram[34][15]=1;ram[34][16]=0;ram[34][17]=1;ram[34][18]=1;ram[34][19]=0;ram[34][20]=0;ram[34][21]=1;ram[34][22]=1;ram[34][23]=0;ram[34][24]=1;ram[34][25]=1;ram[34][26]=1;ram[34][27]=1;ram[34][28]=1;ram[34][29]=1;ram[34][30]=1;ram[34][31]=1;ram[34][32]=1;ram[34][33]=1;ram[34][34]=1;ram[34][35]=0;ram[34][36]=1;ram[34][37]=0;ram[34][38]=0;ram[34][39]=0;ram[34][40]=1;ram[34][41]=0;ram[34][42]=1;ram[34][43]=0;ram[34][44]=1;ram[34][45]=0;ram[34][46]=1;ram[34][47]=0;ram[34][48]=1;ram[34][49]=0;ram[34][50]=1;ram[34][51]=1;ram[34][52]=1;ram[34][53]=1;ram[34][54]=1;ram[34][55]=1;ram[34][56]=1;ram[34][57]=0;ram[34][58]=1;ram[34][59]=0;ram[34][60]=1;ram[34][61]=1;ram[34][62]=0;ram[34][63]=0;ram[34][64]=0;ram[34][65]=1;ram[34][66]=1;ram[34][67]=1;ram[34][68]=1;ram[34][69]=0;ram[34][70]=0;ram[34][71]=0;ram[34][72]=1;ram[34][73]=0;ram[34][74]=1;ram[34][75]=1;ram[34][76]=1;ram[34][77]=1;ram[34][78]=0;ram[34][79]=0;ram[34][80]=0;ram[34][81]=1;ram[34][82]=1;ram[34][83]=0;ram[34][84]=1;ram[34][85]=1;ram[34][86]=0;ram[34][87]=0;ram[34][88]=1;ram[34][89]=1;ram[34][90]=1;ram[34][91]=0;ram[34][92]=1;ram[34][93]=1;ram[34][94]=1;ram[34][95]=0;ram[34][96]=1;ram[34][97]=1;ram[34][98]=0;ram[34][99]=1;ram[34][100]=0;ram[34][101]=1;ram[34][102]=0;ram[34][103]=1;ram[34][104]=1;ram[34][105]=1;ram[34][106]=1;ram[34][107]=1;ram[34][108]=1;ram[34][109]=1;ram[34][110]=1;ram[34][111]=0;ram[34][112]=1;ram[34][113]=1;ram[34][114]=1;ram[34][115]=1;ram[34][116]=0;ram[34][117]=1;ram[34][118]=1;ram[34][119]=0;ram[34][120]=0;ram[34][121]=0;ram[34][122]=1;ram[34][123]=1;ram[34][124]=1;ram[34][125]=1;ram[34][126]=1;ram[34][127]=1;ram[34][128]=0;ram[34][129]=0;ram[34][130]=1;ram[34][131]=1;ram[34][132]=1;ram[34][133]=0;ram[34][134]=0;ram[34][135]=1;ram[34][136]=1;
        ram[35][0]=0;ram[35][1]=1;ram[35][2]=1;ram[35][3]=1;ram[35][4]=1;ram[35][5]=1;ram[35][6]=0;ram[35][7]=1;ram[35][8]=0;ram[35][9]=1;ram[35][10]=1;ram[35][11]=1;ram[35][12]=0;ram[35][13]=1;ram[35][14]=1;ram[35][15]=1;ram[35][16]=1;ram[35][17]=0;ram[35][18]=1;ram[35][19]=1;ram[35][20]=1;ram[35][21]=1;ram[35][22]=1;ram[35][23]=1;ram[35][24]=1;ram[35][25]=1;ram[35][26]=1;ram[35][27]=1;ram[35][28]=1;ram[35][29]=1;ram[35][30]=0;ram[35][31]=1;ram[35][32]=1;ram[35][33]=0;ram[35][34]=1;ram[35][35]=1;ram[35][36]=1;ram[35][37]=0;ram[35][38]=1;ram[35][39]=1;ram[35][40]=0;ram[35][41]=0;ram[35][42]=1;ram[35][43]=0;ram[35][44]=0;ram[35][45]=1;ram[35][46]=1;ram[35][47]=1;ram[35][48]=1;ram[35][49]=1;ram[35][50]=1;ram[35][51]=0;ram[35][52]=0;ram[35][53]=1;ram[35][54]=0;ram[35][55]=0;ram[35][56]=1;ram[35][57]=1;ram[35][58]=0;ram[35][59]=0;ram[35][60]=1;ram[35][61]=1;ram[35][62]=1;ram[35][63]=1;ram[35][64]=0;ram[35][65]=0;ram[35][66]=1;ram[35][67]=1;ram[35][68]=1;ram[35][69]=1;ram[35][70]=0;ram[35][71]=1;ram[35][72]=1;ram[35][73]=0;ram[35][74]=0;ram[35][75]=1;ram[35][76]=1;ram[35][77]=1;ram[35][78]=1;ram[35][79]=1;ram[35][80]=1;ram[35][81]=0;ram[35][82]=0;ram[35][83]=1;ram[35][84]=1;ram[35][85]=1;ram[35][86]=1;ram[35][87]=1;ram[35][88]=1;ram[35][89]=0;ram[35][90]=1;ram[35][91]=1;ram[35][92]=0;ram[35][93]=1;ram[35][94]=1;ram[35][95]=1;ram[35][96]=0;ram[35][97]=1;ram[35][98]=1;ram[35][99]=1;ram[35][100]=1;ram[35][101]=1;ram[35][102]=1;ram[35][103]=1;ram[35][104]=1;ram[35][105]=0;ram[35][106]=0;ram[35][107]=1;ram[35][108]=0;ram[35][109]=0;ram[35][110]=1;ram[35][111]=1;ram[35][112]=0;ram[35][113]=1;ram[35][114]=1;ram[35][115]=0;ram[35][116]=1;ram[35][117]=1;ram[35][118]=1;ram[35][119]=0;ram[35][120]=1;ram[35][121]=1;ram[35][122]=1;ram[35][123]=1;ram[35][124]=1;ram[35][125]=1;ram[35][126]=1;ram[35][127]=1;ram[35][128]=1;ram[35][129]=1;ram[35][130]=0;ram[35][131]=0;ram[35][132]=0;ram[35][133]=0;ram[35][134]=1;ram[35][135]=1;ram[35][136]=0;
        ram[36][0]=1;ram[36][1]=1;ram[36][2]=1;ram[36][3]=0;ram[36][4]=1;ram[36][5]=1;ram[36][6]=1;ram[36][7]=0;ram[36][8]=1;ram[36][9]=1;ram[36][10]=1;ram[36][11]=1;ram[36][12]=1;ram[36][13]=1;ram[36][14]=1;ram[36][15]=1;ram[36][16]=1;ram[36][17]=1;ram[36][18]=0;ram[36][19]=0;ram[36][20]=0;ram[36][21]=1;ram[36][22]=0;ram[36][23]=1;ram[36][24]=0;ram[36][25]=0;ram[36][26]=1;ram[36][27]=1;ram[36][28]=1;ram[36][29]=0;ram[36][30]=1;ram[36][31]=0;ram[36][32]=1;ram[36][33]=1;ram[36][34]=0;ram[36][35]=1;ram[36][36]=1;ram[36][37]=0;ram[36][38]=1;ram[36][39]=1;ram[36][40]=1;ram[36][41]=1;ram[36][42]=1;ram[36][43]=0;ram[36][44]=0;ram[36][45]=1;ram[36][46]=1;ram[36][47]=1;ram[36][48]=1;ram[36][49]=1;ram[36][50]=0;ram[36][51]=1;ram[36][52]=1;ram[36][53]=1;ram[36][54]=1;ram[36][55]=0;ram[36][56]=1;ram[36][57]=0;ram[36][58]=1;ram[36][59]=1;ram[36][60]=0;ram[36][61]=1;ram[36][62]=0;ram[36][63]=1;ram[36][64]=1;ram[36][65]=1;ram[36][66]=1;ram[36][67]=0;ram[36][68]=0;ram[36][69]=1;ram[36][70]=1;ram[36][71]=1;ram[36][72]=0;ram[36][73]=0;ram[36][74]=1;ram[36][75]=0;ram[36][76]=1;ram[36][77]=0;ram[36][78]=0;ram[36][79]=1;ram[36][80]=0;ram[36][81]=1;ram[36][82]=1;ram[36][83]=1;ram[36][84]=1;ram[36][85]=1;ram[36][86]=1;ram[36][87]=0;ram[36][88]=1;ram[36][89]=0;ram[36][90]=1;ram[36][91]=1;ram[36][92]=1;ram[36][93]=1;ram[36][94]=1;ram[36][95]=1;ram[36][96]=0;ram[36][97]=1;ram[36][98]=0;ram[36][99]=1;ram[36][100]=0;ram[36][101]=1;ram[36][102]=0;ram[36][103]=1;ram[36][104]=1;ram[36][105]=1;ram[36][106]=1;ram[36][107]=1;ram[36][108]=0;ram[36][109]=0;ram[36][110]=0;ram[36][111]=1;ram[36][112]=1;ram[36][113]=0;ram[36][114]=1;ram[36][115]=1;ram[36][116]=1;ram[36][117]=1;ram[36][118]=1;ram[36][119]=0;ram[36][120]=1;ram[36][121]=1;ram[36][122]=1;ram[36][123]=1;ram[36][124]=1;ram[36][125]=1;ram[36][126]=1;ram[36][127]=1;ram[36][128]=1;ram[36][129]=1;ram[36][130]=1;ram[36][131]=1;ram[36][132]=1;ram[36][133]=1;ram[36][134]=1;ram[36][135]=1;ram[36][136]=1;
        ram[37][0]=1;ram[37][1]=1;ram[37][2]=1;ram[37][3]=0;ram[37][4]=1;ram[37][5]=1;ram[37][6]=0;ram[37][7]=1;ram[37][8]=1;ram[37][9]=1;ram[37][10]=0;ram[37][11]=0;ram[37][12]=0;ram[37][13]=1;ram[37][14]=0;ram[37][15]=0;ram[37][16]=1;ram[37][17]=0;ram[37][18]=0;ram[37][19]=1;ram[37][20]=0;ram[37][21]=1;ram[37][22]=1;ram[37][23]=1;ram[37][24]=0;ram[37][25]=1;ram[37][26]=1;ram[37][27]=1;ram[37][28]=1;ram[37][29]=0;ram[37][30]=1;ram[37][31]=0;ram[37][32]=1;ram[37][33]=1;ram[37][34]=1;ram[37][35]=1;ram[37][36]=0;ram[37][37]=0;ram[37][38]=1;ram[37][39]=1;ram[37][40]=1;ram[37][41]=0;ram[37][42]=0;ram[37][43]=1;ram[37][44]=1;ram[37][45]=0;ram[37][46]=1;ram[37][47]=1;ram[37][48]=1;ram[37][49]=1;ram[37][50]=1;ram[37][51]=1;ram[37][52]=0;ram[37][53]=1;ram[37][54]=1;ram[37][55]=1;ram[37][56]=1;ram[37][57]=1;ram[37][58]=1;ram[37][59]=1;ram[37][60]=1;ram[37][61]=0;ram[37][62]=1;ram[37][63]=1;ram[37][64]=1;ram[37][65]=1;ram[37][66]=1;ram[37][67]=1;ram[37][68]=1;ram[37][69]=1;ram[37][70]=1;ram[37][71]=1;ram[37][72]=1;ram[37][73]=1;ram[37][74]=1;ram[37][75]=0;ram[37][76]=0;ram[37][77]=0;ram[37][78]=1;ram[37][79]=0;ram[37][80]=1;ram[37][81]=0;ram[37][82]=0;ram[37][83]=0;ram[37][84]=1;ram[37][85]=0;ram[37][86]=1;ram[37][87]=0;ram[37][88]=1;ram[37][89]=0;ram[37][90]=1;ram[37][91]=1;ram[37][92]=1;ram[37][93]=1;ram[37][94]=1;ram[37][95]=1;ram[37][96]=1;ram[37][97]=1;ram[37][98]=0;ram[37][99]=1;ram[37][100]=1;ram[37][101]=0;ram[37][102]=1;ram[37][103]=0;ram[37][104]=0;ram[37][105]=1;ram[37][106]=1;ram[37][107]=0;ram[37][108]=1;ram[37][109]=0;ram[37][110]=0;ram[37][111]=1;ram[37][112]=1;ram[37][113]=1;ram[37][114]=1;ram[37][115]=0;ram[37][116]=0;ram[37][117]=1;ram[37][118]=1;ram[37][119]=1;ram[37][120]=1;ram[37][121]=1;ram[37][122]=1;ram[37][123]=0;ram[37][124]=1;ram[37][125]=1;ram[37][126]=1;ram[37][127]=1;ram[37][128]=1;ram[37][129]=1;ram[37][130]=1;ram[37][131]=1;ram[37][132]=1;ram[37][133]=1;ram[37][134]=1;ram[37][135]=0;ram[37][136]=1;
        ram[38][0]=0;ram[38][1]=1;ram[38][2]=0;ram[38][3]=0;ram[38][4]=1;ram[38][5]=0;ram[38][6]=1;ram[38][7]=0;ram[38][8]=1;ram[38][9]=1;ram[38][10]=1;ram[38][11]=1;ram[38][12]=1;ram[38][13]=0;ram[38][14]=1;ram[38][15]=1;ram[38][16]=1;ram[38][17]=0;ram[38][18]=1;ram[38][19]=0;ram[38][20]=1;ram[38][21]=1;ram[38][22]=1;ram[38][23]=0;ram[38][24]=0;ram[38][25]=1;ram[38][26]=1;ram[38][27]=1;ram[38][28]=1;ram[38][29]=1;ram[38][30]=0;ram[38][31]=1;ram[38][32]=0;ram[38][33]=0;ram[38][34]=1;ram[38][35]=1;ram[38][36]=1;ram[38][37]=1;ram[38][38]=1;ram[38][39]=1;ram[38][40]=1;ram[38][41]=1;ram[38][42]=1;ram[38][43]=1;ram[38][44]=0;ram[38][45]=0;ram[38][46]=1;ram[38][47]=0;ram[38][48]=1;ram[38][49]=1;ram[38][50]=1;ram[38][51]=1;ram[38][52]=1;ram[38][53]=0;ram[38][54]=0;ram[38][55]=0;ram[38][56]=1;ram[38][57]=1;ram[38][58]=1;ram[38][59]=1;ram[38][60]=1;ram[38][61]=1;ram[38][62]=1;ram[38][63]=1;ram[38][64]=1;ram[38][65]=1;ram[38][66]=0;ram[38][67]=0;ram[38][68]=1;ram[38][69]=0;ram[38][70]=0;ram[38][71]=1;ram[38][72]=1;ram[38][73]=1;ram[38][74]=0;ram[38][75]=0;ram[38][76]=0;ram[38][77]=1;ram[38][78]=1;ram[38][79]=1;ram[38][80]=1;ram[38][81]=1;ram[38][82]=0;ram[38][83]=1;ram[38][84]=1;ram[38][85]=1;ram[38][86]=0;ram[38][87]=0;ram[38][88]=1;ram[38][89]=1;ram[38][90]=1;ram[38][91]=1;ram[38][92]=1;ram[38][93]=1;ram[38][94]=1;ram[38][95]=0;ram[38][96]=1;ram[38][97]=0;ram[38][98]=1;ram[38][99]=0;ram[38][100]=0;ram[38][101]=0;ram[38][102]=1;ram[38][103]=1;ram[38][104]=1;ram[38][105]=0;ram[38][106]=0;ram[38][107]=1;ram[38][108]=0;ram[38][109]=1;ram[38][110]=0;ram[38][111]=0;ram[38][112]=0;ram[38][113]=1;ram[38][114]=0;ram[38][115]=1;ram[38][116]=1;ram[38][117]=0;ram[38][118]=1;ram[38][119]=1;ram[38][120]=1;ram[38][121]=1;ram[38][122]=0;ram[38][123]=1;ram[38][124]=1;ram[38][125]=1;ram[38][126]=1;ram[38][127]=1;ram[38][128]=0;ram[38][129]=0;ram[38][130]=1;ram[38][131]=1;ram[38][132]=0;ram[38][133]=1;ram[38][134]=0;ram[38][135]=1;ram[38][136]=1;
        ram[39][0]=1;ram[39][1]=0;ram[39][2]=0;ram[39][3]=1;ram[39][4]=1;ram[39][5]=1;ram[39][6]=0;ram[39][7]=1;ram[39][8]=1;ram[39][9]=1;ram[39][10]=1;ram[39][11]=1;ram[39][12]=1;ram[39][13]=0;ram[39][14]=1;ram[39][15]=1;ram[39][16]=1;ram[39][17]=0;ram[39][18]=1;ram[39][19]=1;ram[39][20]=1;ram[39][21]=1;ram[39][22]=1;ram[39][23]=1;ram[39][24]=1;ram[39][25]=1;ram[39][26]=1;ram[39][27]=1;ram[39][28]=0;ram[39][29]=1;ram[39][30]=1;ram[39][31]=1;ram[39][32]=0;ram[39][33]=1;ram[39][34]=1;ram[39][35]=1;ram[39][36]=1;ram[39][37]=1;ram[39][38]=1;ram[39][39]=0;ram[39][40]=1;ram[39][41]=1;ram[39][42]=1;ram[39][43]=1;ram[39][44]=1;ram[39][45]=0;ram[39][46]=0;ram[39][47]=1;ram[39][48]=1;ram[39][49]=1;ram[39][50]=1;ram[39][51]=1;ram[39][52]=1;ram[39][53]=1;ram[39][54]=1;ram[39][55]=1;ram[39][56]=0;ram[39][57]=1;ram[39][58]=1;ram[39][59]=0;ram[39][60]=1;ram[39][61]=0;ram[39][62]=0;ram[39][63]=1;ram[39][64]=1;ram[39][65]=0;ram[39][66]=1;ram[39][67]=1;ram[39][68]=1;ram[39][69]=1;ram[39][70]=1;ram[39][71]=0;ram[39][72]=1;ram[39][73]=1;ram[39][74]=0;ram[39][75]=0;ram[39][76]=0;ram[39][77]=1;ram[39][78]=1;ram[39][79]=0;ram[39][80]=1;ram[39][81]=1;ram[39][82]=1;ram[39][83]=1;ram[39][84]=1;ram[39][85]=1;ram[39][86]=0;ram[39][87]=1;ram[39][88]=1;ram[39][89]=1;ram[39][90]=1;ram[39][91]=1;ram[39][92]=1;ram[39][93]=0;ram[39][94]=0;ram[39][95]=1;ram[39][96]=1;ram[39][97]=1;ram[39][98]=1;ram[39][99]=0;ram[39][100]=1;ram[39][101]=1;ram[39][102]=1;ram[39][103]=1;ram[39][104]=1;ram[39][105]=1;ram[39][106]=1;ram[39][107]=0;ram[39][108]=1;ram[39][109]=1;ram[39][110]=1;ram[39][111]=1;ram[39][112]=1;ram[39][113]=0;ram[39][114]=0;ram[39][115]=1;ram[39][116]=1;ram[39][117]=1;ram[39][118]=0;ram[39][119]=1;ram[39][120]=1;ram[39][121]=1;ram[39][122]=1;ram[39][123]=0;ram[39][124]=1;ram[39][125]=1;ram[39][126]=0;ram[39][127]=1;ram[39][128]=1;ram[39][129]=1;ram[39][130]=1;ram[39][131]=0;ram[39][132]=1;ram[39][133]=1;ram[39][134]=0;ram[39][135]=1;ram[39][136]=0;
        ram[40][0]=1;ram[40][1]=0;ram[40][2]=1;ram[40][3]=1;ram[40][4]=0;ram[40][5]=1;ram[40][6]=1;ram[40][7]=1;ram[40][8]=0;ram[40][9]=1;ram[40][10]=0;ram[40][11]=1;ram[40][12]=0;ram[40][13]=0;ram[40][14]=1;ram[40][15]=0;ram[40][16]=1;ram[40][17]=1;ram[40][18]=0;ram[40][19]=0;ram[40][20]=1;ram[40][21]=0;ram[40][22]=1;ram[40][23]=1;ram[40][24]=0;ram[40][25]=0;ram[40][26]=1;ram[40][27]=1;ram[40][28]=1;ram[40][29]=1;ram[40][30]=1;ram[40][31]=0;ram[40][32]=1;ram[40][33]=1;ram[40][34]=1;ram[40][35]=1;ram[40][36]=0;ram[40][37]=1;ram[40][38]=0;ram[40][39]=1;ram[40][40]=0;ram[40][41]=0;ram[40][42]=1;ram[40][43]=0;ram[40][44]=1;ram[40][45]=1;ram[40][46]=0;ram[40][47]=1;ram[40][48]=0;ram[40][49]=1;ram[40][50]=1;ram[40][51]=1;ram[40][52]=1;ram[40][53]=1;ram[40][54]=0;ram[40][55]=0;ram[40][56]=1;ram[40][57]=1;ram[40][58]=0;ram[40][59]=1;ram[40][60]=0;ram[40][61]=1;ram[40][62]=1;ram[40][63]=1;ram[40][64]=1;ram[40][65]=1;ram[40][66]=0;ram[40][67]=1;ram[40][68]=1;ram[40][69]=1;ram[40][70]=0;ram[40][71]=1;ram[40][72]=1;ram[40][73]=0;ram[40][74]=1;ram[40][75]=1;ram[40][76]=1;ram[40][77]=1;ram[40][78]=0;ram[40][79]=0;ram[40][80]=1;ram[40][81]=1;ram[40][82]=0;ram[40][83]=0;ram[40][84]=1;ram[40][85]=0;ram[40][86]=0;ram[40][87]=1;ram[40][88]=0;ram[40][89]=1;ram[40][90]=0;ram[40][91]=0;ram[40][92]=0;ram[40][93]=1;ram[40][94]=1;ram[40][95]=0;ram[40][96]=0;ram[40][97]=1;ram[40][98]=1;ram[40][99]=1;ram[40][100]=0;ram[40][101]=1;ram[40][102]=1;ram[40][103]=1;ram[40][104]=0;ram[40][105]=1;ram[40][106]=1;ram[40][107]=1;ram[40][108]=1;ram[40][109]=0;ram[40][110]=0;ram[40][111]=1;ram[40][112]=0;ram[40][113]=1;ram[40][114]=1;ram[40][115]=1;ram[40][116]=0;ram[40][117]=1;ram[40][118]=1;ram[40][119]=0;ram[40][120]=1;ram[40][121]=0;ram[40][122]=0;ram[40][123]=1;ram[40][124]=1;ram[40][125]=1;ram[40][126]=1;ram[40][127]=1;ram[40][128]=1;ram[40][129]=1;ram[40][130]=1;ram[40][131]=1;ram[40][132]=1;ram[40][133]=0;ram[40][134]=1;ram[40][135]=0;ram[40][136]=0;
        ram[41][0]=1;ram[41][1]=1;ram[41][2]=0;ram[41][3]=1;ram[41][4]=0;ram[41][5]=1;ram[41][6]=1;ram[41][7]=0;ram[41][8]=1;ram[41][9]=0;ram[41][10]=1;ram[41][11]=1;ram[41][12]=0;ram[41][13]=1;ram[41][14]=1;ram[41][15]=0;ram[41][16]=1;ram[41][17]=0;ram[41][18]=1;ram[41][19]=1;ram[41][20]=1;ram[41][21]=1;ram[41][22]=1;ram[41][23]=1;ram[41][24]=1;ram[41][25]=1;ram[41][26]=1;ram[41][27]=1;ram[41][28]=1;ram[41][29]=0;ram[41][30]=0;ram[41][31]=1;ram[41][32]=0;ram[41][33]=0;ram[41][34]=1;ram[41][35]=1;ram[41][36]=0;ram[41][37]=1;ram[41][38]=1;ram[41][39]=0;ram[41][40]=1;ram[41][41]=0;ram[41][42]=0;ram[41][43]=1;ram[41][44]=1;ram[41][45]=0;ram[41][46]=1;ram[41][47]=1;ram[41][48]=1;ram[41][49]=1;ram[41][50]=0;ram[41][51]=1;ram[41][52]=0;ram[41][53]=1;ram[41][54]=0;ram[41][55]=1;ram[41][56]=1;ram[41][57]=1;ram[41][58]=1;ram[41][59]=1;ram[41][60]=1;ram[41][61]=0;ram[41][62]=1;ram[41][63]=0;ram[41][64]=1;ram[41][65]=1;ram[41][66]=1;ram[41][67]=1;ram[41][68]=1;ram[41][69]=1;ram[41][70]=1;ram[41][71]=1;ram[41][72]=1;ram[41][73]=1;ram[41][74]=1;ram[41][75]=1;ram[41][76]=1;ram[41][77]=1;ram[41][78]=1;ram[41][79]=1;ram[41][80]=0;ram[41][81]=0;ram[41][82]=1;ram[41][83]=1;ram[41][84]=0;ram[41][85]=0;ram[41][86]=1;ram[41][87]=1;ram[41][88]=0;ram[41][89]=1;ram[41][90]=0;ram[41][91]=1;ram[41][92]=1;ram[41][93]=1;ram[41][94]=1;ram[41][95]=1;ram[41][96]=0;ram[41][97]=1;ram[41][98]=0;ram[41][99]=0;ram[41][100]=1;ram[41][101]=0;ram[41][102]=1;ram[41][103]=1;ram[41][104]=0;ram[41][105]=0;ram[41][106]=1;ram[41][107]=1;ram[41][108]=1;ram[41][109]=1;ram[41][110]=0;ram[41][111]=1;ram[41][112]=1;ram[41][113]=0;ram[41][114]=1;ram[41][115]=1;ram[41][116]=0;ram[41][117]=0;ram[41][118]=1;ram[41][119]=0;ram[41][120]=1;ram[41][121]=0;ram[41][122]=1;ram[41][123]=1;ram[41][124]=0;ram[41][125]=0;ram[41][126]=1;ram[41][127]=1;ram[41][128]=1;ram[41][129]=1;ram[41][130]=0;ram[41][131]=1;ram[41][132]=0;ram[41][133]=0;ram[41][134]=1;ram[41][135]=0;ram[41][136]=0;
        ram[42][0]=1;ram[42][1]=1;ram[42][2]=0;ram[42][3]=0;ram[42][4]=1;ram[42][5]=0;ram[42][6]=1;ram[42][7]=1;ram[42][8]=1;ram[42][9]=1;ram[42][10]=0;ram[42][11]=1;ram[42][12]=1;ram[42][13]=0;ram[42][14]=0;ram[42][15]=1;ram[42][16]=1;ram[42][17]=1;ram[42][18]=1;ram[42][19]=1;ram[42][20]=0;ram[42][21]=0;ram[42][22]=0;ram[42][23]=1;ram[42][24]=0;ram[42][25]=1;ram[42][26]=1;ram[42][27]=0;ram[42][28]=0;ram[42][29]=1;ram[42][30]=1;ram[42][31]=0;ram[42][32]=0;ram[42][33]=1;ram[42][34]=0;ram[42][35]=1;ram[42][36]=0;ram[42][37]=1;ram[42][38]=0;ram[42][39]=1;ram[42][40]=1;ram[42][41]=1;ram[42][42]=0;ram[42][43]=1;ram[42][44]=0;ram[42][45]=0;ram[42][46]=0;ram[42][47]=1;ram[42][48]=1;ram[42][49]=0;ram[42][50]=1;ram[42][51]=1;ram[42][52]=1;ram[42][53]=1;ram[42][54]=1;ram[42][55]=0;ram[42][56]=0;ram[42][57]=1;ram[42][58]=0;ram[42][59]=1;ram[42][60]=1;ram[42][61]=0;ram[42][62]=1;ram[42][63]=0;ram[42][64]=1;ram[42][65]=1;ram[42][66]=1;ram[42][67]=0;ram[42][68]=0;ram[42][69]=1;ram[42][70]=0;ram[42][71]=1;ram[42][72]=1;ram[42][73]=1;ram[42][74]=1;ram[42][75]=1;ram[42][76]=1;ram[42][77]=0;ram[42][78]=1;ram[42][79]=1;ram[42][80]=1;ram[42][81]=1;ram[42][82]=1;ram[42][83]=1;ram[42][84]=1;ram[42][85]=1;ram[42][86]=1;ram[42][87]=1;ram[42][88]=1;ram[42][89]=0;ram[42][90]=1;ram[42][91]=0;ram[42][92]=1;ram[42][93]=1;ram[42][94]=0;ram[42][95]=0;ram[42][96]=0;ram[42][97]=1;ram[42][98]=0;ram[42][99]=1;ram[42][100]=1;ram[42][101]=0;ram[42][102]=0;ram[42][103]=1;ram[42][104]=0;ram[42][105]=1;ram[42][106]=0;ram[42][107]=0;ram[42][108]=0;ram[42][109]=1;ram[42][110]=0;ram[42][111]=0;ram[42][112]=1;ram[42][113]=1;ram[42][114]=1;ram[42][115]=1;ram[42][116]=0;ram[42][117]=1;ram[42][118]=0;ram[42][119]=1;ram[42][120]=0;ram[42][121]=0;ram[42][122]=0;ram[42][123]=1;ram[42][124]=1;ram[42][125]=1;ram[42][126]=1;ram[42][127]=0;ram[42][128]=0;ram[42][129]=0;ram[42][130]=1;ram[42][131]=0;ram[42][132]=0;ram[42][133]=1;ram[42][134]=1;ram[42][135]=0;ram[42][136]=0;
        ram[43][0]=1;ram[43][1]=1;ram[43][2]=1;ram[43][3]=0;ram[43][4]=1;ram[43][5]=1;ram[43][6]=1;ram[43][7]=1;ram[43][8]=0;ram[43][9]=0;ram[43][10]=1;ram[43][11]=0;ram[43][12]=0;ram[43][13]=1;ram[43][14]=0;ram[43][15]=1;ram[43][16]=1;ram[43][17]=0;ram[43][18]=1;ram[43][19]=0;ram[43][20]=1;ram[43][21]=1;ram[43][22]=0;ram[43][23]=1;ram[43][24]=0;ram[43][25]=1;ram[43][26]=1;ram[43][27]=1;ram[43][28]=0;ram[43][29]=1;ram[43][30]=1;ram[43][31]=0;ram[43][32]=1;ram[43][33]=1;ram[43][34]=1;ram[43][35]=0;ram[43][36]=0;ram[43][37]=1;ram[43][38]=0;ram[43][39]=1;ram[43][40]=0;ram[43][41]=0;ram[43][42]=1;ram[43][43]=0;ram[43][44]=0;ram[43][45]=1;ram[43][46]=1;ram[43][47]=1;ram[43][48]=1;ram[43][49]=0;ram[43][50]=0;ram[43][51]=0;ram[43][52]=0;ram[43][53]=1;ram[43][54]=1;ram[43][55]=0;ram[43][56]=1;ram[43][57]=0;ram[43][58]=1;ram[43][59]=0;ram[43][60]=1;ram[43][61]=1;ram[43][62]=1;ram[43][63]=0;ram[43][64]=1;ram[43][65]=1;ram[43][66]=1;ram[43][67]=0;ram[43][68]=1;ram[43][69]=1;ram[43][70]=0;ram[43][71]=1;ram[43][72]=0;ram[43][73]=1;ram[43][74]=1;ram[43][75]=0;ram[43][76]=0;ram[43][77]=1;ram[43][78]=1;ram[43][79]=1;ram[43][80]=1;ram[43][81]=1;ram[43][82]=1;ram[43][83]=1;ram[43][84]=1;ram[43][85]=1;ram[43][86]=1;ram[43][87]=1;ram[43][88]=0;ram[43][89]=0;ram[43][90]=1;ram[43][91]=1;ram[43][92]=1;ram[43][93]=1;ram[43][94]=0;ram[43][95]=0;ram[43][96]=0;ram[43][97]=1;ram[43][98]=1;ram[43][99]=1;ram[43][100]=1;ram[43][101]=1;ram[43][102]=0;ram[43][103]=1;ram[43][104]=0;ram[43][105]=0;ram[43][106]=1;ram[43][107]=0;ram[43][108]=1;ram[43][109]=0;ram[43][110]=1;ram[43][111]=1;ram[43][112]=1;ram[43][113]=0;ram[43][114]=1;ram[43][115]=1;ram[43][116]=1;ram[43][117]=1;ram[43][118]=0;ram[43][119]=1;ram[43][120]=0;ram[43][121]=1;ram[43][122]=0;ram[43][123]=1;ram[43][124]=0;ram[43][125]=1;ram[43][126]=0;ram[43][127]=0;ram[43][128]=1;ram[43][129]=1;ram[43][130]=1;ram[43][131]=0;ram[43][132]=1;ram[43][133]=1;ram[43][134]=0;ram[43][135]=1;ram[43][136]=0;
        ram[44][0]=1;ram[44][1]=1;ram[44][2]=0;ram[44][3]=1;ram[44][4]=1;ram[44][5]=1;ram[44][6]=1;ram[44][7]=0;ram[44][8]=1;ram[44][9]=0;ram[44][10]=1;ram[44][11]=1;ram[44][12]=1;ram[44][13]=0;ram[44][14]=1;ram[44][15]=1;ram[44][16]=1;ram[44][17]=1;ram[44][18]=1;ram[44][19]=1;ram[44][20]=1;ram[44][21]=1;ram[44][22]=0;ram[44][23]=0;ram[44][24]=1;ram[44][25]=1;ram[44][26]=1;ram[44][27]=1;ram[44][28]=1;ram[44][29]=1;ram[44][30]=0;ram[44][31]=1;ram[44][32]=1;ram[44][33]=0;ram[44][34]=0;ram[44][35]=1;ram[44][36]=1;ram[44][37]=1;ram[44][38]=1;ram[44][39]=0;ram[44][40]=1;ram[44][41]=1;ram[44][42]=1;ram[44][43]=0;ram[44][44]=0;ram[44][45]=1;ram[44][46]=1;ram[44][47]=1;ram[44][48]=1;ram[44][49]=1;ram[44][50]=1;ram[44][51]=1;ram[44][52]=1;ram[44][53]=0;ram[44][54]=1;ram[44][55]=1;ram[44][56]=0;ram[44][57]=0;ram[44][58]=1;ram[44][59]=1;ram[44][60]=0;ram[44][61]=0;ram[44][62]=1;ram[44][63]=1;ram[44][64]=1;ram[44][65]=1;ram[44][66]=1;ram[44][67]=0;ram[44][68]=1;ram[44][69]=1;ram[44][70]=1;ram[44][71]=1;ram[44][72]=0;ram[44][73]=1;ram[44][74]=0;ram[44][75]=1;ram[44][76]=0;ram[44][77]=1;ram[44][78]=0;ram[44][79]=1;ram[44][80]=0;ram[44][81]=1;ram[44][82]=0;ram[44][83]=1;ram[44][84]=1;ram[44][85]=0;ram[44][86]=0;ram[44][87]=0;ram[44][88]=0;ram[44][89]=0;ram[44][90]=0;ram[44][91]=1;ram[44][92]=1;ram[44][93]=1;ram[44][94]=0;ram[44][95]=0;ram[44][96]=1;ram[44][97]=0;ram[44][98]=1;ram[44][99]=0;ram[44][100]=0;ram[44][101]=1;ram[44][102]=0;ram[44][103]=1;ram[44][104]=1;ram[44][105]=1;ram[44][106]=0;ram[44][107]=0;ram[44][108]=0;ram[44][109]=1;ram[44][110]=1;ram[44][111]=1;ram[44][112]=1;ram[44][113]=1;ram[44][114]=1;ram[44][115]=0;ram[44][116]=0;ram[44][117]=0;ram[44][118]=1;ram[44][119]=1;ram[44][120]=1;ram[44][121]=1;ram[44][122]=1;ram[44][123]=1;ram[44][124]=1;ram[44][125]=1;ram[44][126]=1;ram[44][127]=0;ram[44][128]=1;ram[44][129]=0;ram[44][130]=1;ram[44][131]=0;ram[44][132]=1;ram[44][133]=1;ram[44][134]=1;ram[44][135]=1;ram[44][136]=0;
        ram[45][0]=0;ram[45][1]=1;ram[45][2]=1;ram[45][3]=0;ram[45][4]=1;ram[45][5]=1;ram[45][6]=1;ram[45][7]=1;ram[45][8]=1;ram[45][9]=1;ram[45][10]=0;ram[45][11]=1;ram[45][12]=1;ram[45][13]=1;ram[45][14]=1;ram[45][15]=1;ram[45][16]=1;ram[45][17]=0;ram[45][18]=1;ram[45][19]=1;ram[45][20]=1;ram[45][21]=1;ram[45][22]=1;ram[45][23]=0;ram[45][24]=1;ram[45][25]=1;ram[45][26]=1;ram[45][27]=1;ram[45][28]=0;ram[45][29]=1;ram[45][30]=1;ram[45][31]=1;ram[45][32]=0;ram[45][33]=1;ram[45][34]=1;ram[45][35]=0;ram[45][36]=1;ram[45][37]=1;ram[45][38]=0;ram[45][39]=0;ram[45][40]=1;ram[45][41]=1;ram[45][42]=1;ram[45][43]=1;ram[45][44]=0;ram[45][45]=0;ram[45][46]=1;ram[45][47]=0;ram[45][48]=1;ram[45][49]=1;ram[45][50]=1;ram[45][51]=1;ram[45][52]=1;ram[45][53]=0;ram[45][54]=1;ram[45][55]=0;ram[45][56]=1;ram[45][57]=1;ram[45][58]=1;ram[45][59]=1;ram[45][60]=0;ram[45][61]=1;ram[45][62]=1;ram[45][63]=1;ram[45][64]=1;ram[45][65]=1;ram[45][66]=1;ram[45][67]=0;ram[45][68]=1;ram[45][69]=0;ram[45][70]=1;ram[45][71]=1;ram[45][72]=1;ram[45][73]=0;ram[45][74]=0;ram[45][75]=1;ram[45][76]=0;ram[45][77]=1;ram[45][78]=0;ram[45][79]=0;ram[45][80]=1;ram[45][81]=0;ram[45][82]=1;ram[45][83]=0;ram[45][84]=1;ram[45][85]=0;ram[45][86]=0;ram[45][87]=1;ram[45][88]=0;ram[45][89]=1;ram[45][90]=0;ram[45][91]=0;ram[45][92]=1;ram[45][93]=0;ram[45][94]=0;ram[45][95]=1;ram[45][96]=1;ram[45][97]=0;ram[45][98]=0;ram[45][99]=0;ram[45][100]=1;ram[45][101]=0;ram[45][102]=1;ram[45][103]=0;ram[45][104]=0;ram[45][105]=0;ram[45][106]=1;ram[45][107]=0;ram[45][108]=0;ram[45][109]=0;ram[45][110]=1;ram[45][111]=1;ram[45][112]=0;ram[45][113]=1;ram[45][114]=0;ram[45][115]=0;ram[45][116]=0;ram[45][117]=1;ram[45][118]=1;ram[45][119]=0;ram[45][120]=1;ram[45][121]=0;ram[45][122]=1;ram[45][123]=1;ram[45][124]=1;ram[45][125]=0;ram[45][126]=0;ram[45][127]=1;ram[45][128]=0;ram[45][129]=1;ram[45][130]=1;ram[45][131]=1;ram[45][132]=1;ram[45][133]=1;ram[45][134]=0;ram[45][135]=0;ram[45][136]=0;
        ram[46][0]=1;ram[46][1]=0;ram[46][2]=1;ram[46][3]=1;ram[46][4]=0;ram[46][5]=1;ram[46][6]=1;ram[46][7]=0;ram[46][8]=0;ram[46][9]=0;ram[46][10]=1;ram[46][11]=1;ram[46][12]=1;ram[46][13]=0;ram[46][14]=1;ram[46][15]=0;ram[46][16]=1;ram[46][17]=1;ram[46][18]=1;ram[46][19]=0;ram[46][20]=0;ram[46][21]=0;ram[46][22]=0;ram[46][23]=1;ram[46][24]=1;ram[46][25]=0;ram[46][26]=1;ram[46][27]=1;ram[46][28]=0;ram[46][29]=1;ram[46][30]=0;ram[46][31]=1;ram[46][32]=1;ram[46][33]=1;ram[46][34]=1;ram[46][35]=0;ram[46][36]=1;ram[46][37]=1;ram[46][38]=0;ram[46][39]=0;ram[46][40]=1;ram[46][41]=1;ram[46][42]=0;ram[46][43]=1;ram[46][44]=1;ram[46][45]=1;ram[46][46]=1;ram[46][47]=1;ram[46][48]=0;ram[46][49]=1;ram[46][50]=1;ram[46][51]=0;ram[46][52]=0;ram[46][53]=1;ram[46][54]=1;ram[46][55]=0;ram[46][56]=1;ram[46][57]=1;ram[46][58]=1;ram[46][59]=1;ram[46][60]=1;ram[46][61]=1;ram[46][62]=1;ram[46][63]=1;ram[46][64]=1;ram[46][65]=0;ram[46][66]=0;ram[46][67]=1;ram[46][68]=1;ram[46][69]=0;ram[46][70]=1;ram[46][71]=1;ram[46][72]=0;ram[46][73]=0;ram[46][74]=0;ram[46][75]=1;ram[46][76]=0;ram[46][77]=1;ram[46][78]=1;ram[46][79]=1;ram[46][80]=0;ram[46][81]=1;ram[46][82]=0;ram[46][83]=1;ram[46][84]=0;ram[46][85]=1;ram[46][86]=1;ram[46][87]=1;ram[46][88]=0;ram[46][89]=1;ram[46][90]=1;ram[46][91]=0;ram[46][92]=0;ram[46][93]=0;ram[46][94]=1;ram[46][95]=0;ram[46][96]=1;ram[46][97]=0;ram[46][98]=1;ram[46][99]=0;ram[46][100]=0;ram[46][101]=1;ram[46][102]=1;ram[46][103]=1;ram[46][104]=1;ram[46][105]=1;ram[46][106]=0;ram[46][107]=0;ram[46][108]=0;ram[46][109]=0;ram[46][110]=0;ram[46][111]=0;ram[46][112]=0;ram[46][113]=0;ram[46][114]=0;ram[46][115]=1;ram[46][116]=1;ram[46][117]=1;ram[46][118]=1;ram[46][119]=0;ram[46][120]=1;ram[46][121]=0;ram[46][122]=1;ram[46][123]=1;ram[46][124]=0;ram[46][125]=1;ram[46][126]=0;ram[46][127]=0;ram[46][128]=0;ram[46][129]=1;ram[46][130]=1;ram[46][131]=1;ram[46][132]=0;ram[46][133]=1;ram[46][134]=0;ram[46][135]=1;ram[46][136]=1;
        ram[47][0]=0;ram[47][1]=1;ram[47][2]=0;ram[47][3]=1;ram[47][4]=0;ram[47][5]=0;ram[47][6]=1;ram[47][7]=1;ram[47][8]=1;ram[47][9]=1;ram[47][10]=0;ram[47][11]=1;ram[47][12]=0;ram[47][13]=1;ram[47][14]=1;ram[47][15]=1;ram[47][16]=0;ram[47][17]=1;ram[47][18]=1;ram[47][19]=1;ram[47][20]=1;ram[47][21]=0;ram[47][22]=0;ram[47][23]=1;ram[47][24]=0;ram[47][25]=0;ram[47][26]=1;ram[47][27]=0;ram[47][28]=1;ram[47][29]=0;ram[47][30]=1;ram[47][31]=1;ram[47][32]=0;ram[47][33]=1;ram[47][34]=0;ram[47][35]=1;ram[47][36]=1;ram[47][37]=0;ram[47][38]=0;ram[47][39]=1;ram[47][40]=0;ram[47][41]=1;ram[47][42]=1;ram[47][43]=1;ram[47][44]=1;ram[47][45]=0;ram[47][46]=1;ram[47][47]=1;ram[47][48]=1;ram[47][49]=0;ram[47][50]=1;ram[47][51]=0;ram[47][52]=1;ram[47][53]=0;ram[47][54]=1;ram[47][55]=1;ram[47][56]=1;ram[47][57]=1;ram[47][58]=0;ram[47][59]=1;ram[47][60]=0;ram[47][61]=0;ram[47][62]=0;ram[47][63]=1;ram[47][64]=1;ram[47][65]=1;ram[47][66]=1;ram[47][67]=1;ram[47][68]=1;ram[47][69]=1;ram[47][70]=1;ram[47][71]=1;ram[47][72]=1;ram[47][73]=1;ram[47][74]=1;ram[47][75]=1;ram[47][76]=1;ram[47][77]=0;ram[47][78]=1;ram[47][79]=1;ram[47][80]=0;ram[47][81]=1;ram[47][82]=0;ram[47][83]=0;ram[47][84]=1;ram[47][85]=1;ram[47][86]=1;ram[47][87]=1;ram[47][88]=0;ram[47][89]=1;ram[47][90]=1;ram[47][91]=0;ram[47][92]=1;ram[47][93]=0;ram[47][94]=1;ram[47][95]=1;ram[47][96]=0;ram[47][97]=1;ram[47][98]=0;ram[47][99]=0;ram[47][100]=1;ram[47][101]=1;ram[47][102]=0;ram[47][103]=1;ram[47][104]=1;ram[47][105]=1;ram[47][106]=0;ram[47][107]=1;ram[47][108]=1;ram[47][109]=1;ram[47][110]=1;ram[47][111]=1;ram[47][112]=0;ram[47][113]=0;ram[47][114]=1;ram[47][115]=1;ram[47][116]=1;ram[47][117]=0;ram[47][118]=1;ram[47][119]=1;ram[47][120]=1;ram[47][121]=1;ram[47][122]=1;ram[47][123]=1;ram[47][124]=0;ram[47][125]=1;ram[47][126]=1;ram[47][127]=1;ram[47][128]=0;ram[47][129]=1;ram[47][130]=1;ram[47][131]=1;ram[47][132]=1;ram[47][133]=0;ram[47][134]=1;ram[47][135]=1;ram[47][136]=0;
        ram[48][0]=1;ram[48][1]=1;ram[48][2]=1;ram[48][3]=0;ram[48][4]=1;ram[48][5]=0;ram[48][6]=1;ram[48][7]=0;ram[48][8]=1;ram[48][9]=0;ram[48][10]=1;ram[48][11]=1;ram[48][12]=0;ram[48][13]=0;ram[48][14]=1;ram[48][15]=0;ram[48][16]=1;ram[48][17]=1;ram[48][18]=1;ram[48][19]=1;ram[48][20]=1;ram[48][21]=0;ram[48][22]=1;ram[48][23]=0;ram[48][24]=1;ram[48][25]=1;ram[48][26]=1;ram[48][27]=1;ram[48][28]=1;ram[48][29]=1;ram[48][30]=1;ram[48][31]=1;ram[48][32]=1;ram[48][33]=1;ram[48][34]=1;ram[48][35]=1;ram[48][36]=1;ram[48][37]=0;ram[48][38]=0;ram[48][39]=0;ram[48][40]=0;ram[48][41]=1;ram[48][42]=1;ram[48][43]=1;ram[48][44]=1;ram[48][45]=0;ram[48][46]=1;ram[48][47]=0;ram[48][48]=1;ram[48][49]=0;ram[48][50]=1;ram[48][51]=1;ram[48][52]=1;ram[48][53]=1;ram[48][54]=0;ram[48][55]=1;ram[48][56]=0;ram[48][57]=1;ram[48][58]=0;ram[48][59]=0;ram[48][60]=0;ram[48][61]=1;ram[48][62]=1;ram[48][63]=1;ram[48][64]=1;ram[48][65]=0;ram[48][66]=0;ram[48][67]=1;ram[48][68]=1;ram[48][69]=0;ram[48][70]=0;ram[48][71]=1;ram[48][72]=1;ram[48][73]=1;ram[48][74]=1;ram[48][75]=1;ram[48][76]=0;ram[48][77]=1;ram[48][78]=1;ram[48][79]=1;ram[48][80]=1;ram[48][81]=1;ram[48][82]=1;ram[48][83]=0;ram[48][84]=1;ram[48][85]=1;ram[48][86]=0;ram[48][87]=1;ram[48][88]=1;ram[48][89]=1;ram[48][90]=0;ram[48][91]=0;ram[48][92]=1;ram[48][93]=0;ram[48][94]=1;ram[48][95]=1;ram[48][96]=1;ram[48][97]=1;ram[48][98]=1;ram[48][99]=0;ram[48][100]=1;ram[48][101]=0;ram[48][102]=1;ram[48][103]=1;ram[48][104]=1;ram[48][105]=1;ram[48][106]=1;ram[48][107]=0;ram[48][108]=1;ram[48][109]=0;ram[48][110]=0;ram[48][111]=1;ram[48][112]=1;ram[48][113]=1;ram[48][114]=1;ram[48][115]=1;ram[48][116]=1;ram[48][117]=1;ram[48][118]=1;ram[48][119]=0;ram[48][120]=1;ram[48][121]=0;ram[48][122]=1;ram[48][123]=0;ram[48][124]=0;ram[48][125]=0;ram[48][126]=1;ram[48][127]=1;ram[48][128]=1;ram[48][129]=1;ram[48][130]=0;ram[48][131]=1;ram[48][132]=1;ram[48][133]=1;ram[48][134]=0;ram[48][135]=0;ram[48][136]=0;
        ram[49][0]=0;ram[49][1]=0;ram[49][2]=1;ram[49][3]=1;ram[49][4]=1;ram[49][5]=1;ram[49][6]=1;ram[49][7]=1;ram[49][8]=1;ram[49][9]=1;ram[49][10]=1;ram[49][11]=0;ram[49][12]=0;ram[49][13]=1;ram[49][14]=0;ram[49][15]=0;ram[49][16]=1;ram[49][17]=0;ram[49][18]=1;ram[49][19]=1;ram[49][20]=1;ram[49][21]=1;ram[49][22]=0;ram[49][23]=1;ram[49][24]=1;ram[49][25]=1;ram[49][26]=0;ram[49][27]=1;ram[49][28]=0;ram[49][29]=1;ram[49][30]=1;ram[49][31]=1;ram[49][32]=0;ram[49][33]=0;ram[49][34]=0;ram[49][35]=1;ram[49][36]=1;ram[49][37]=0;ram[49][38]=1;ram[49][39]=0;ram[49][40]=1;ram[49][41]=1;ram[49][42]=0;ram[49][43]=1;ram[49][44]=1;ram[49][45]=1;ram[49][46]=0;ram[49][47]=1;ram[49][48]=1;ram[49][49]=0;ram[49][50]=1;ram[49][51]=0;ram[49][52]=1;ram[49][53]=1;ram[49][54]=1;ram[49][55]=0;ram[49][56]=1;ram[49][57]=0;ram[49][58]=1;ram[49][59]=0;ram[49][60]=0;ram[49][61]=1;ram[49][62]=0;ram[49][63]=1;ram[49][64]=1;ram[49][65]=1;ram[49][66]=0;ram[49][67]=0;ram[49][68]=1;ram[49][69]=1;ram[49][70]=1;ram[49][71]=0;ram[49][72]=1;ram[49][73]=1;ram[49][74]=0;ram[49][75]=1;ram[49][76]=0;ram[49][77]=1;ram[49][78]=1;ram[49][79]=0;ram[49][80]=1;ram[49][81]=1;ram[49][82]=1;ram[49][83]=1;ram[49][84]=1;ram[49][85]=1;ram[49][86]=0;ram[49][87]=0;ram[49][88]=0;ram[49][89]=1;ram[49][90]=0;ram[49][91]=0;ram[49][92]=0;ram[49][93]=1;ram[49][94]=1;ram[49][95]=0;ram[49][96]=0;ram[49][97]=0;ram[49][98]=0;ram[49][99]=0;ram[49][100]=0;ram[49][101]=1;ram[49][102]=1;ram[49][103]=1;ram[49][104]=0;ram[49][105]=1;ram[49][106]=0;ram[49][107]=1;ram[49][108]=1;ram[49][109]=1;ram[49][110]=1;ram[49][111]=0;ram[49][112]=1;ram[49][113]=1;ram[49][114]=1;ram[49][115]=0;ram[49][116]=0;ram[49][117]=1;ram[49][118]=0;ram[49][119]=0;ram[49][120]=1;ram[49][121]=0;ram[49][122]=0;ram[49][123]=0;ram[49][124]=1;ram[49][125]=1;ram[49][126]=1;ram[49][127]=1;ram[49][128]=1;ram[49][129]=0;ram[49][130]=1;ram[49][131]=1;ram[49][132]=1;ram[49][133]=1;ram[49][134]=0;ram[49][135]=1;ram[49][136]=1;
        ram[50][0]=1;ram[50][1]=0;ram[50][2]=1;ram[50][3]=1;ram[50][4]=1;ram[50][5]=1;ram[50][6]=0;ram[50][7]=0;ram[50][8]=1;ram[50][9]=1;ram[50][10]=1;ram[50][11]=1;ram[50][12]=0;ram[50][13]=0;ram[50][14]=0;ram[50][15]=1;ram[50][16]=1;ram[50][17]=0;ram[50][18]=0;ram[50][19]=1;ram[50][20]=0;ram[50][21]=0;ram[50][22]=1;ram[50][23]=1;ram[50][24]=1;ram[50][25]=1;ram[50][26]=1;ram[50][27]=1;ram[50][28]=0;ram[50][29]=1;ram[50][30]=1;ram[50][31]=1;ram[50][32]=1;ram[50][33]=1;ram[50][34]=0;ram[50][35]=0;ram[50][36]=1;ram[50][37]=1;ram[50][38]=0;ram[50][39]=1;ram[50][40]=0;ram[50][41]=1;ram[50][42]=0;ram[50][43]=0;ram[50][44]=0;ram[50][45]=1;ram[50][46]=0;ram[50][47]=1;ram[50][48]=1;ram[50][49]=0;ram[50][50]=1;ram[50][51]=1;ram[50][52]=0;ram[50][53]=1;ram[50][54]=1;ram[50][55]=1;ram[50][56]=1;ram[50][57]=0;ram[50][58]=1;ram[50][59]=0;ram[50][60]=1;ram[50][61]=1;ram[50][62]=1;ram[50][63]=1;ram[50][64]=0;ram[50][65]=1;ram[50][66]=0;ram[50][67]=0;ram[50][68]=1;ram[50][69]=0;ram[50][70]=1;ram[50][71]=1;ram[50][72]=0;ram[50][73]=0;ram[50][74]=0;ram[50][75]=1;ram[50][76]=0;ram[50][77]=1;ram[50][78]=0;ram[50][79]=0;ram[50][80]=0;ram[50][81]=0;ram[50][82]=0;ram[50][83]=0;ram[50][84]=1;ram[50][85]=1;ram[50][86]=0;ram[50][87]=0;ram[50][88]=1;ram[50][89]=1;ram[50][90]=0;ram[50][91]=1;ram[50][92]=0;ram[50][93]=1;ram[50][94]=1;ram[50][95]=1;ram[50][96]=0;ram[50][97]=1;ram[50][98]=1;ram[50][99]=0;ram[50][100]=1;ram[50][101]=1;ram[50][102]=0;ram[50][103]=1;ram[50][104]=1;ram[50][105]=1;ram[50][106]=0;ram[50][107]=1;ram[50][108]=1;ram[50][109]=1;ram[50][110]=1;ram[50][111]=1;ram[50][112]=1;ram[50][113]=1;ram[50][114]=1;ram[50][115]=1;ram[50][116]=0;ram[50][117]=1;ram[50][118]=1;ram[50][119]=1;ram[50][120]=1;ram[50][121]=0;ram[50][122]=0;ram[50][123]=1;ram[50][124]=0;ram[50][125]=1;ram[50][126]=1;ram[50][127]=1;ram[50][128]=1;ram[50][129]=1;ram[50][130]=0;ram[50][131]=1;ram[50][132]=1;ram[50][133]=1;ram[50][134]=0;ram[50][135]=1;ram[50][136]=1;
        ram[51][0]=1;ram[51][1]=1;ram[51][2]=1;ram[51][3]=0;ram[51][4]=1;ram[51][5]=1;ram[51][6]=0;ram[51][7]=1;ram[51][8]=0;ram[51][9]=0;ram[51][10]=1;ram[51][11]=0;ram[51][12]=0;ram[51][13]=1;ram[51][14]=0;ram[51][15]=0;ram[51][16]=1;ram[51][17]=1;ram[51][18]=1;ram[51][19]=0;ram[51][20]=1;ram[51][21]=1;ram[51][22]=1;ram[51][23]=1;ram[51][24]=1;ram[51][25]=0;ram[51][26]=1;ram[51][27]=1;ram[51][28]=1;ram[51][29]=0;ram[51][30]=0;ram[51][31]=0;ram[51][32]=0;ram[51][33]=0;ram[51][34]=0;ram[51][35]=0;ram[51][36]=1;ram[51][37]=0;ram[51][38]=0;ram[51][39]=1;ram[51][40]=1;ram[51][41]=1;ram[51][42]=1;ram[51][43]=1;ram[51][44]=1;ram[51][45]=1;ram[51][46]=1;ram[51][47]=0;ram[51][48]=0;ram[51][49]=0;ram[51][50]=1;ram[51][51]=0;ram[51][52]=0;ram[51][53]=1;ram[51][54]=1;ram[51][55]=1;ram[51][56]=1;ram[51][57]=1;ram[51][58]=0;ram[51][59]=0;ram[51][60]=1;ram[51][61]=1;ram[51][62]=1;ram[51][63]=1;ram[51][64]=0;ram[51][65]=1;ram[51][66]=0;ram[51][67]=1;ram[51][68]=1;ram[51][69]=0;ram[51][70]=1;ram[51][71]=1;ram[51][72]=0;ram[51][73]=1;ram[51][74]=0;ram[51][75]=1;ram[51][76]=0;ram[51][77]=1;ram[51][78]=1;ram[51][79]=1;ram[51][80]=0;ram[51][81]=1;ram[51][82]=0;ram[51][83]=0;ram[51][84]=1;ram[51][85]=1;ram[51][86]=0;ram[51][87]=0;ram[51][88]=1;ram[51][89]=1;ram[51][90]=1;ram[51][91]=1;ram[51][92]=1;ram[51][93]=0;ram[51][94]=0;ram[51][95]=1;ram[51][96]=1;ram[51][97]=1;ram[51][98]=1;ram[51][99]=1;ram[51][100]=1;ram[51][101]=0;ram[51][102]=1;ram[51][103]=0;ram[51][104]=0;ram[51][105]=0;ram[51][106]=1;ram[51][107]=0;ram[51][108]=1;ram[51][109]=1;ram[51][110]=1;ram[51][111]=0;ram[51][112]=1;ram[51][113]=1;ram[51][114]=1;ram[51][115]=1;ram[51][116]=0;ram[51][117]=1;ram[51][118]=1;ram[51][119]=0;ram[51][120]=1;ram[51][121]=1;ram[51][122]=0;ram[51][123]=1;ram[51][124]=1;ram[51][125]=1;ram[51][126]=0;ram[51][127]=0;ram[51][128]=1;ram[51][129]=1;ram[51][130]=1;ram[51][131]=0;ram[51][132]=0;ram[51][133]=1;ram[51][134]=1;ram[51][135]=1;ram[51][136]=1;
        ram[52][0]=1;ram[52][1]=0;ram[52][2]=1;ram[52][3]=0;ram[52][4]=0;ram[52][5]=1;ram[52][6]=0;ram[52][7]=0;ram[52][8]=0;ram[52][9]=1;ram[52][10]=1;ram[52][11]=1;ram[52][12]=1;ram[52][13]=0;ram[52][14]=1;ram[52][15]=1;ram[52][16]=0;ram[52][17]=0;ram[52][18]=1;ram[52][19]=0;ram[52][20]=0;ram[52][21]=1;ram[52][22]=1;ram[52][23]=1;ram[52][24]=0;ram[52][25]=0;ram[52][26]=1;ram[52][27]=0;ram[52][28]=1;ram[52][29]=0;ram[52][30]=0;ram[52][31]=1;ram[52][32]=1;ram[52][33]=1;ram[52][34]=0;ram[52][35]=1;ram[52][36]=0;ram[52][37]=0;ram[52][38]=0;ram[52][39]=1;ram[52][40]=1;ram[52][41]=1;ram[52][42]=1;ram[52][43]=1;ram[52][44]=1;ram[52][45]=1;ram[52][46]=0;ram[52][47]=0;ram[52][48]=1;ram[52][49]=0;ram[52][50]=1;ram[52][51]=0;ram[52][52]=0;ram[52][53]=0;ram[52][54]=0;ram[52][55]=1;ram[52][56]=1;ram[52][57]=1;ram[52][58]=1;ram[52][59]=1;ram[52][60]=1;ram[52][61]=1;ram[52][62]=1;ram[52][63]=0;ram[52][64]=1;ram[52][65]=1;ram[52][66]=0;ram[52][67]=0;ram[52][68]=1;ram[52][69]=0;ram[52][70]=0;ram[52][71]=0;ram[52][72]=1;ram[52][73]=0;ram[52][74]=1;ram[52][75]=0;ram[52][76]=1;ram[52][77]=0;ram[52][78]=0;ram[52][79]=0;ram[52][80]=0;ram[52][81]=0;ram[52][82]=1;ram[52][83]=1;ram[52][84]=1;ram[52][85]=1;ram[52][86]=0;ram[52][87]=1;ram[52][88]=0;ram[52][89]=0;ram[52][90]=1;ram[52][91]=1;ram[52][92]=0;ram[52][93]=1;ram[52][94]=1;ram[52][95]=1;ram[52][96]=1;ram[52][97]=0;ram[52][98]=0;ram[52][99]=1;ram[52][100]=0;ram[52][101]=0;ram[52][102]=1;ram[52][103]=1;ram[52][104]=0;ram[52][105]=1;ram[52][106]=1;ram[52][107]=0;ram[52][108]=1;ram[52][109]=1;ram[52][110]=0;ram[52][111]=1;ram[52][112]=0;ram[52][113]=0;ram[52][114]=1;ram[52][115]=1;ram[52][116]=0;ram[52][117]=1;ram[52][118]=0;ram[52][119]=1;ram[52][120]=1;ram[52][121]=1;ram[52][122]=1;ram[52][123]=1;ram[52][124]=1;ram[52][125]=1;ram[52][126]=0;ram[52][127]=1;ram[52][128]=1;ram[52][129]=1;ram[52][130]=1;ram[52][131]=1;ram[52][132]=1;ram[52][133]=1;ram[52][134]=1;ram[52][135]=1;ram[52][136]=1;
        ram[53][0]=1;ram[53][1]=1;ram[53][2]=0;ram[53][3]=1;ram[53][4]=1;ram[53][5]=0;ram[53][6]=1;ram[53][7]=0;ram[53][8]=1;ram[53][9]=1;ram[53][10]=1;ram[53][11]=1;ram[53][12]=1;ram[53][13]=1;ram[53][14]=1;ram[53][15]=1;ram[53][16]=1;ram[53][17]=1;ram[53][18]=1;ram[53][19]=1;ram[53][20]=1;ram[53][21]=1;ram[53][22]=1;ram[53][23]=0;ram[53][24]=1;ram[53][25]=0;ram[53][26]=1;ram[53][27]=0;ram[53][28]=1;ram[53][29]=1;ram[53][30]=1;ram[53][31]=1;ram[53][32]=1;ram[53][33]=1;ram[53][34]=1;ram[53][35]=0;ram[53][36]=0;ram[53][37]=0;ram[53][38]=0;ram[53][39]=1;ram[53][40]=1;ram[53][41]=1;ram[53][42]=0;ram[53][43]=1;ram[53][44]=1;ram[53][45]=0;ram[53][46]=1;ram[53][47]=0;ram[53][48]=1;ram[53][49]=1;ram[53][50]=1;ram[53][51]=0;ram[53][52]=0;ram[53][53]=1;ram[53][54]=1;ram[53][55]=1;ram[53][56]=0;ram[53][57]=0;ram[53][58]=1;ram[53][59]=1;ram[53][60]=1;ram[53][61]=1;ram[53][62]=0;ram[53][63]=1;ram[53][64]=1;ram[53][65]=1;ram[53][66]=0;ram[53][67]=1;ram[53][68]=0;ram[53][69]=1;ram[53][70]=1;ram[53][71]=0;ram[53][72]=0;ram[53][73]=0;ram[53][74]=1;ram[53][75]=1;ram[53][76]=1;ram[53][77]=1;ram[53][78]=1;ram[53][79]=1;ram[53][80]=1;ram[53][81]=1;ram[53][82]=1;ram[53][83]=0;ram[53][84]=0;ram[53][85]=1;ram[53][86]=1;ram[53][87]=0;ram[53][88]=1;ram[53][89]=0;ram[53][90]=1;ram[53][91]=1;ram[53][92]=1;ram[53][93]=0;ram[53][94]=0;ram[53][95]=0;ram[53][96]=0;ram[53][97]=1;ram[53][98]=1;ram[53][99]=0;ram[53][100]=1;ram[53][101]=1;ram[53][102]=1;ram[53][103]=1;ram[53][104]=1;ram[53][105]=0;ram[53][106]=1;ram[53][107]=1;ram[53][108]=1;ram[53][109]=1;ram[53][110]=0;ram[53][111]=1;ram[53][112]=1;ram[53][113]=1;ram[53][114]=1;ram[53][115]=1;ram[53][116]=1;ram[53][117]=1;ram[53][118]=1;ram[53][119]=1;ram[53][120]=1;ram[53][121]=1;ram[53][122]=1;ram[53][123]=0;ram[53][124]=1;ram[53][125]=1;ram[53][126]=1;ram[53][127]=1;ram[53][128]=0;ram[53][129]=1;ram[53][130]=0;ram[53][131]=1;ram[53][132]=1;ram[53][133]=0;ram[53][134]=0;ram[53][135]=1;ram[53][136]=1;
        ram[54][0]=0;ram[54][1]=1;ram[54][2]=1;ram[54][3]=0;ram[54][4]=1;ram[54][5]=0;ram[54][6]=0;ram[54][7]=1;ram[54][8]=1;ram[54][9]=1;ram[54][10]=0;ram[54][11]=1;ram[54][12]=0;ram[54][13]=0;ram[54][14]=1;ram[54][15]=0;ram[54][16]=1;ram[54][17]=0;ram[54][18]=1;ram[54][19]=1;ram[54][20]=0;ram[54][21]=1;ram[54][22]=0;ram[54][23]=1;ram[54][24]=1;ram[54][25]=1;ram[54][26]=1;ram[54][27]=0;ram[54][28]=1;ram[54][29]=1;ram[54][30]=0;ram[54][31]=1;ram[54][32]=0;ram[54][33]=1;ram[54][34]=1;ram[54][35]=1;ram[54][36]=0;ram[54][37]=0;ram[54][38]=1;ram[54][39]=1;ram[54][40]=1;ram[54][41]=1;ram[54][42]=1;ram[54][43]=1;ram[54][44]=1;ram[54][45]=1;ram[54][46]=0;ram[54][47]=1;ram[54][48]=1;ram[54][49]=0;ram[54][50]=1;ram[54][51]=0;ram[54][52]=0;ram[54][53]=1;ram[54][54]=1;ram[54][55]=1;ram[54][56]=1;ram[54][57]=1;ram[54][58]=1;ram[54][59]=0;ram[54][60]=1;ram[54][61]=1;ram[54][62]=0;ram[54][63]=1;ram[54][64]=1;ram[54][65]=1;ram[54][66]=1;ram[54][67]=0;ram[54][68]=1;ram[54][69]=1;ram[54][70]=0;ram[54][71]=0;ram[54][72]=1;ram[54][73]=1;ram[54][74]=1;ram[54][75]=0;ram[54][76]=1;ram[54][77]=1;ram[54][78]=1;ram[54][79]=1;ram[54][80]=1;ram[54][81]=1;ram[54][82]=1;ram[54][83]=1;ram[54][84]=0;ram[54][85]=1;ram[54][86]=1;ram[54][87]=1;ram[54][88]=0;ram[54][89]=1;ram[54][90]=1;ram[54][91]=1;ram[54][92]=1;ram[54][93]=0;ram[54][94]=1;ram[54][95]=0;ram[54][96]=0;ram[54][97]=1;ram[54][98]=1;ram[54][99]=0;ram[54][100]=1;ram[54][101]=0;ram[54][102]=1;ram[54][103]=0;ram[54][104]=1;ram[54][105]=1;ram[54][106]=0;ram[54][107]=0;ram[54][108]=1;ram[54][109]=1;ram[54][110]=1;ram[54][111]=0;ram[54][112]=1;ram[54][113]=0;ram[54][114]=0;ram[54][115]=1;ram[54][116]=1;ram[54][117]=1;ram[54][118]=1;ram[54][119]=0;ram[54][120]=1;ram[54][121]=0;ram[54][122]=1;ram[54][123]=1;ram[54][124]=0;ram[54][125]=1;ram[54][126]=1;ram[54][127]=1;ram[54][128]=0;ram[54][129]=1;ram[54][130]=0;ram[54][131]=0;ram[54][132]=0;ram[54][133]=0;ram[54][134]=1;ram[54][135]=0;ram[54][136]=0;
        ram[55][0]=0;ram[55][1]=0;ram[55][2]=0;ram[55][3]=1;ram[55][4]=1;ram[55][5]=1;ram[55][6]=1;ram[55][7]=1;ram[55][8]=0;ram[55][9]=1;ram[55][10]=1;ram[55][11]=1;ram[55][12]=1;ram[55][13]=1;ram[55][14]=1;ram[55][15]=0;ram[55][16]=1;ram[55][17]=1;ram[55][18]=1;ram[55][19]=1;ram[55][20]=1;ram[55][21]=0;ram[55][22]=0;ram[55][23]=1;ram[55][24]=0;ram[55][25]=1;ram[55][26]=1;ram[55][27]=1;ram[55][28]=1;ram[55][29]=1;ram[55][30]=0;ram[55][31]=1;ram[55][32]=1;ram[55][33]=1;ram[55][34]=0;ram[55][35]=1;ram[55][36]=1;ram[55][37]=1;ram[55][38]=0;ram[55][39]=1;ram[55][40]=1;ram[55][41]=1;ram[55][42]=1;ram[55][43]=1;ram[55][44]=1;ram[55][45]=0;ram[55][46]=1;ram[55][47]=1;ram[55][48]=1;ram[55][49]=1;ram[55][50]=1;ram[55][51]=0;ram[55][52]=1;ram[55][53]=1;ram[55][54]=1;ram[55][55]=1;ram[55][56]=1;ram[55][57]=0;ram[55][58]=1;ram[55][59]=0;ram[55][60]=1;ram[55][61]=0;ram[55][62]=1;ram[55][63]=1;ram[55][64]=0;ram[55][65]=1;ram[55][66]=0;ram[55][67]=0;ram[55][68]=1;ram[55][69]=1;ram[55][70]=1;ram[55][71]=1;ram[55][72]=0;ram[55][73]=0;ram[55][74]=0;ram[55][75]=0;ram[55][76]=1;ram[55][77]=1;ram[55][78]=1;ram[55][79]=1;ram[55][80]=1;ram[55][81]=0;ram[55][82]=0;ram[55][83]=0;ram[55][84]=1;ram[55][85]=1;ram[55][86]=0;ram[55][87]=1;ram[55][88]=0;ram[55][89]=1;ram[55][90]=0;ram[55][91]=0;ram[55][92]=1;ram[55][93]=1;ram[55][94]=1;ram[55][95]=1;ram[55][96]=1;ram[55][97]=1;ram[55][98]=1;ram[55][99]=1;ram[55][100]=1;ram[55][101]=1;ram[55][102]=1;ram[55][103]=1;ram[55][104]=0;ram[55][105]=0;ram[55][106]=0;ram[55][107]=0;ram[55][108]=1;ram[55][109]=0;ram[55][110]=1;ram[55][111]=1;ram[55][112]=1;ram[55][113]=1;ram[55][114]=1;ram[55][115]=1;ram[55][116]=1;ram[55][117]=1;ram[55][118]=1;ram[55][119]=0;ram[55][120]=1;ram[55][121]=1;ram[55][122]=1;ram[55][123]=1;ram[55][124]=1;ram[55][125]=1;ram[55][126]=1;ram[55][127]=1;ram[55][128]=1;ram[55][129]=1;ram[55][130]=1;ram[55][131]=1;ram[55][132]=1;ram[55][133]=0;ram[55][134]=1;ram[55][135]=1;ram[55][136]=1;
        ram[56][0]=1;ram[56][1]=1;ram[56][2]=0;ram[56][3]=0;ram[56][4]=1;ram[56][5]=0;ram[56][6]=1;ram[56][7]=1;ram[56][8]=1;ram[56][9]=1;ram[56][10]=1;ram[56][11]=1;ram[56][12]=1;ram[56][13]=0;ram[56][14]=0;ram[56][15]=1;ram[56][16]=1;ram[56][17]=1;ram[56][18]=1;ram[56][19]=1;ram[56][20]=0;ram[56][21]=1;ram[56][22]=0;ram[56][23]=1;ram[56][24]=1;ram[56][25]=1;ram[56][26]=0;ram[56][27]=0;ram[56][28]=0;ram[56][29]=1;ram[56][30]=1;ram[56][31]=1;ram[56][32]=0;ram[56][33]=1;ram[56][34]=1;ram[56][35]=0;ram[56][36]=1;ram[56][37]=1;ram[56][38]=1;ram[56][39]=1;ram[56][40]=1;ram[56][41]=0;ram[56][42]=0;ram[56][43]=1;ram[56][44]=1;ram[56][45]=1;ram[56][46]=1;ram[56][47]=1;ram[56][48]=1;ram[56][49]=0;ram[56][50]=1;ram[56][51]=1;ram[56][52]=1;ram[56][53]=1;ram[56][54]=1;ram[56][55]=1;ram[56][56]=1;ram[56][57]=1;ram[56][58]=1;ram[56][59]=1;ram[56][60]=1;ram[56][61]=1;ram[56][62]=0;ram[56][63]=1;ram[56][64]=1;ram[56][65]=0;ram[56][66]=1;ram[56][67]=0;ram[56][68]=0;ram[56][69]=1;ram[56][70]=1;ram[56][71]=1;ram[56][72]=0;ram[56][73]=1;ram[56][74]=1;ram[56][75]=0;ram[56][76]=0;ram[56][77]=0;ram[56][78]=0;ram[56][79]=0;ram[56][80]=0;ram[56][81]=1;ram[56][82]=1;ram[56][83]=1;ram[56][84]=0;ram[56][85]=1;ram[56][86]=1;ram[56][87]=1;ram[56][88]=0;ram[56][89]=0;ram[56][90]=1;ram[56][91]=0;ram[56][92]=0;ram[56][93]=0;ram[56][94]=0;ram[56][95]=1;ram[56][96]=1;ram[56][97]=0;ram[56][98]=1;ram[56][99]=1;ram[56][100]=1;ram[56][101]=1;ram[56][102]=0;ram[56][103]=0;ram[56][104]=0;ram[56][105]=1;ram[56][106]=1;ram[56][107]=1;ram[56][108]=1;ram[56][109]=1;ram[56][110]=1;ram[56][111]=1;ram[56][112]=0;ram[56][113]=1;ram[56][114]=1;ram[56][115]=1;ram[56][116]=1;ram[56][117]=1;ram[56][118]=1;ram[56][119]=1;ram[56][120]=1;ram[56][121]=0;ram[56][122]=0;ram[56][123]=1;ram[56][124]=1;ram[56][125]=1;ram[56][126]=1;ram[56][127]=0;ram[56][128]=1;ram[56][129]=1;ram[56][130]=1;ram[56][131]=0;ram[56][132]=1;ram[56][133]=0;ram[56][134]=1;ram[56][135]=0;ram[56][136]=1;
        ram[57][0]=1;ram[57][1]=1;ram[57][2]=1;ram[57][3]=1;ram[57][4]=1;ram[57][5]=1;ram[57][6]=1;ram[57][7]=1;ram[57][8]=0;ram[57][9]=1;ram[57][10]=0;ram[57][11]=1;ram[57][12]=0;ram[57][13]=1;ram[57][14]=1;ram[57][15]=1;ram[57][16]=0;ram[57][17]=0;ram[57][18]=1;ram[57][19]=1;ram[57][20]=1;ram[57][21]=0;ram[57][22]=1;ram[57][23]=1;ram[57][24]=1;ram[57][25]=0;ram[57][26]=1;ram[57][27]=1;ram[57][28]=1;ram[57][29]=1;ram[57][30]=1;ram[57][31]=1;ram[57][32]=1;ram[57][33]=1;ram[57][34]=0;ram[57][35]=1;ram[57][36]=0;ram[57][37]=0;ram[57][38]=0;ram[57][39]=1;ram[57][40]=1;ram[57][41]=1;ram[57][42]=1;ram[57][43]=0;ram[57][44]=1;ram[57][45]=1;ram[57][46]=1;ram[57][47]=1;ram[57][48]=0;ram[57][49]=1;ram[57][50]=1;ram[57][51]=0;ram[57][52]=0;ram[57][53]=0;ram[57][54]=1;ram[57][55]=1;ram[57][56]=0;ram[57][57]=1;ram[57][58]=0;ram[57][59]=0;ram[57][60]=1;ram[57][61]=0;ram[57][62]=1;ram[57][63]=1;ram[57][64]=0;ram[57][65]=1;ram[57][66]=0;ram[57][67]=0;ram[57][68]=0;ram[57][69]=0;ram[57][70]=0;ram[57][71]=1;ram[57][72]=1;ram[57][73]=1;ram[57][74]=0;ram[57][75]=1;ram[57][76]=0;ram[57][77]=1;ram[57][78]=1;ram[57][79]=1;ram[57][80]=1;ram[57][81]=1;ram[57][82]=1;ram[57][83]=1;ram[57][84]=1;ram[57][85]=1;ram[57][86]=1;ram[57][87]=1;ram[57][88]=1;ram[57][89]=1;ram[57][90]=0;ram[57][91]=1;ram[57][92]=0;ram[57][93]=1;ram[57][94]=1;ram[57][95]=1;ram[57][96]=1;ram[57][97]=0;ram[57][98]=0;ram[57][99]=1;ram[57][100]=0;ram[57][101]=0;ram[57][102]=0;ram[57][103]=1;ram[57][104]=0;ram[57][105]=1;ram[57][106]=0;ram[57][107]=1;ram[57][108]=0;ram[57][109]=1;ram[57][110]=1;ram[57][111]=1;ram[57][112]=0;ram[57][113]=1;ram[57][114]=1;ram[57][115]=0;ram[57][116]=1;ram[57][117]=0;ram[57][118]=0;ram[57][119]=1;ram[57][120]=1;ram[57][121]=0;ram[57][122]=1;ram[57][123]=1;ram[57][124]=1;ram[57][125]=1;ram[57][126]=1;ram[57][127]=0;ram[57][128]=0;ram[57][129]=1;ram[57][130]=0;ram[57][131]=1;ram[57][132]=1;ram[57][133]=1;ram[57][134]=1;ram[57][135]=0;ram[57][136]=0;
        ram[58][0]=1;ram[58][1]=0;ram[58][2]=1;ram[58][3]=0;ram[58][4]=1;ram[58][5]=0;ram[58][6]=0;ram[58][7]=1;ram[58][8]=1;ram[58][9]=1;ram[58][10]=0;ram[58][11]=1;ram[58][12]=1;ram[58][13]=1;ram[58][14]=1;ram[58][15]=1;ram[58][16]=0;ram[58][17]=1;ram[58][18]=0;ram[58][19]=0;ram[58][20]=0;ram[58][21]=1;ram[58][22]=1;ram[58][23]=1;ram[58][24]=1;ram[58][25]=1;ram[58][26]=0;ram[58][27]=1;ram[58][28]=1;ram[58][29]=1;ram[58][30]=1;ram[58][31]=1;ram[58][32]=0;ram[58][33]=1;ram[58][34]=0;ram[58][35]=1;ram[58][36]=1;ram[58][37]=1;ram[58][38]=0;ram[58][39]=1;ram[58][40]=0;ram[58][41]=0;ram[58][42]=1;ram[58][43]=1;ram[58][44]=0;ram[58][45]=1;ram[58][46]=1;ram[58][47]=1;ram[58][48]=0;ram[58][49]=0;ram[58][50]=1;ram[58][51]=0;ram[58][52]=1;ram[58][53]=0;ram[58][54]=1;ram[58][55]=1;ram[58][56]=0;ram[58][57]=1;ram[58][58]=0;ram[58][59]=1;ram[58][60]=0;ram[58][61]=1;ram[58][62]=1;ram[58][63]=0;ram[58][64]=0;ram[58][65]=1;ram[58][66]=1;ram[58][67]=1;ram[58][68]=0;ram[58][69]=1;ram[58][70]=1;ram[58][71]=1;ram[58][72]=1;ram[58][73]=1;ram[58][74]=0;ram[58][75]=0;ram[58][76]=0;ram[58][77]=1;ram[58][78]=1;ram[58][79]=1;ram[58][80]=1;ram[58][81]=1;ram[58][82]=1;ram[58][83]=1;ram[58][84]=0;ram[58][85]=1;ram[58][86]=0;ram[58][87]=1;ram[58][88]=1;ram[58][89]=0;ram[58][90]=1;ram[58][91]=1;ram[58][92]=0;ram[58][93]=0;ram[58][94]=1;ram[58][95]=0;ram[58][96]=0;ram[58][97]=1;ram[58][98]=1;ram[58][99]=0;ram[58][100]=0;ram[58][101]=0;ram[58][102]=1;ram[58][103]=0;ram[58][104]=0;ram[58][105]=0;ram[58][106]=0;ram[58][107]=0;ram[58][108]=0;ram[58][109]=0;ram[58][110]=1;ram[58][111]=1;ram[58][112]=1;ram[58][113]=0;ram[58][114]=1;ram[58][115]=1;ram[58][116]=0;ram[58][117]=1;ram[58][118]=0;ram[58][119]=1;ram[58][120]=1;ram[58][121]=1;ram[58][122]=1;ram[58][123]=0;ram[58][124]=0;ram[58][125]=0;ram[58][126]=0;ram[58][127]=1;ram[58][128]=0;ram[58][129]=1;ram[58][130]=0;ram[58][131]=1;ram[58][132]=0;ram[58][133]=0;ram[58][134]=1;ram[58][135]=1;ram[58][136]=1;
        ram[59][0]=1;ram[59][1]=0;ram[59][2]=1;ram[59][3]=0;ram[59][4]=1;ram[59][5]=1;ram[59][6]=0;ram[59][7]=0;ram[59][8]=0;ram[59][9]=1;ram[59][10]=1;ram[59][11]=1;ram[59][12]=1;ram[59][13]=1;ram[59][14]=1;ram[59][15]=1;ram[59][16]=1;ram[59][17]=0;ram[59][18]=1;ram[59][19]=1;ram[59][20]=1;ram[59][21]=1;ram[59][22]=0;ram[59][23]=1;ram[59][24]=1;ram[59][25]=0;ram[59][26]=1;ram[59][27]=1;ram[59][28]=0;ram[59][29]=1;ram[59][30]=1;ram[59][31]=1;ram[59][32]=1;ram[59][33]=1;ram[59][34]=0;ram[59][35]=0;ram[59][36]=0;ram[59][37]=1;ram[59][38]=1;ram[59][39]=0;ram[59][40]=1;ram[59][41]=0;ram[59][42]=1;ram[59][43]=1;ram[59][44]=1;ram[59][45]=0;ram[59][46]=1;ram[59][47]=1;ram[59][48]=0;ram[59][49]=0;ram[59][50]=0;ram[59][51]=1;ram[59][52]=1;ram[59][53]=0;ram[59][54]=1;ram[59][55]=0;ram[59][56]=0;ram[59][57]=1;ram[59][58]=0;ram[59][59]=1;ram[59][60]=1;ram[59][61]=1;ram[59][62]=0;ram[59][63]=1;ram[59][64]=0;ram[59][65]=1;ram[59][66]=0;ram[59][67]=1;ram[59][68]=1;ram[59][69]=0;ram[59][70]=1;ram[59][71]=1;ram[59][72]=0;ram[59][73]=0;ram[59][74]=1;ram[59][75]=0;ram[59][76]=1;ram[59][77]=1;ram[59][78]=0;ram[59][79]=1;ram[59][80]=0;ram[59][81]=0;ram[59][82]=1;ram[59][83]=1;ram[59][84]=0;ram[59][85]=1;ram[59][86]=1;ram[59][87]=1;ram[59][88]=1;ram[59][89]=0;ram[59][90]=1;ram[59][91]=0;ram[59][92]=0;ram[59][93]=0;ram[59][94]=1;ram[59][95]=1;ram[59][96]=1;ram[59][97]=1;ram[59][98]=1;ram[59][99]=1;ram[59][100]=0;ram[59][101]=0;ram[59][102]=1;ram[59][103]=1;ram[59][104]=0;ram[59][105]=0;ram[59][106]=1;ram[59][107]=0;ram[59][108]=1;ram[59][109]=0;ram[59][110]=0;ram[59][111]=1;ram[59][112]=0;ram[59][113]=0;ram[59][114]=1;ram[59][115]=1;ram[59][116]=0;ram[59][117]=1;ram[59][118]=0;ram[59][119]=1;ram[59][120]=1;ram[59][121]=1;ram[59][122]=1;ram[59][123]=0;ram[59][124]=1;ram[59][125]=0;ram[59][126]=0;ram[59][127]=1;ram[59][128]=1;ram[59][129]=0;ram[59][130]=1;ram[59][131]=0;ram[59][132]=0;ram[59][133]=0;ram[59][134]=0;ram[59][135]=1;ram[59][136]=0;
        ram[60][0]=0;ram[60][1]=1;ram[60][2]=0;ram[60][3]=0;ram[60][4]=1;ram[60][5]=1;ram[60][6]=1;ram[60][7]=1;ram[60][8]=1;ram[60][9]=0;ram[60][10]=0;ram[60][11]=1;ram[60][12]=1;ram[60][13]=1;ram[60][14]=1;ram[60][15]=0;ram[60][16]=0;ram[60][17]=1;ram[60][18]=1;ram[60][19]=1;ram[60][20]=1;ram[60][21]=1;ram[60][22]=0;ram[60][23]=1;ram[60][24]=1;ram[60][25]=1;ram[60][26]=1;ram[60][27]=0;ram[60][28]=1;ram[60][29]=1;ram[60][30]=1;ram[60][31]=1;ram[60][32]=0;ram[60][33]=1;ram[60][34]=1;ram[60][35]=0;ram[60][36]=1;ram[60][37]=1;ram[60][38]=0;ram[60][39]=0;ram[60][40]=1;ram[60][41]=1;ram[60][42]=1;ram[60][43]=0;ram[60][44]=1;ram[60][45]=1;ram[60][46]=1;ram[60][47]=1;ram[60][48]=0;ram[60][49]=0;ram[60][50]=0;ram[60][51]=0;ram[60][52]=0;ram[60][53]=0;ram[60][54]=1;ram[60][55]=1;ram[60][56]=1;ram[60][57]=1;ram[60][58]=1;ram[60][59]=1;ram[60][60]=1;ram[60][61]=1;ram[60][62]=1;ram[60][63]=1;ram[60][64]=1;ram[60][65]=1;ram[60][66]=0;ram[60][67]=1;ram[60][68]=1;ram[60][69]=0;ram[60][70]=0;ram[60][71]=0;ram[60][72]=0;ram[60][73]=1;ram[60][74]=1;ram[60][75]=1;ram[60][76]=0;ram[60][77]=1;ram[60][78]=0;ram[60][79]=1;ram[60][80]=1;ram[60][81]=1;ram[60][82]=1;ram[60][83]=0;ram[60][84]=1;ram[60][85]=1;ram[60][86]=0;ram[60][87]=0;ram[60][88]=0;ram[60][89]=1;ram[60][90]=1;ram[60][91]=0;ram[60][92]=0;ram[60][93]=1;ram[60][94]=1;ram[60][95]=1;ram[60][96]=1;ram[60][97]=0;ram[60][98]=0;ram[60][99]=0;ram[60][100]=1;ram[60][101]=1;ram[60][102]=0;ram[60][103]=1;ram[60][104]=1;ram[60][105]=1;ram[60][106]=1;ram[60][107]=0;ram[60][108]=1;ram[60][109]=1;ram[60][110]=0;ram[60][111]=1;ram[60][112]=1;ram[60][113]=1;ram[60][114]=1;ram[60][115]=1;ram[60][116]=0;ram[60][117]=0;ram[60][118]=1;ram[60][119]=1;ram[60][120]=1;ram[60][121]=1;ram[60][122]=0;ram[60][123]=0;ram[60][124]=1;ram[60][125]=0;ram[60][126]=1;ram[60][127]=0;ram[60][128]=1;ram[60][129]=0;ram[60][130]=1;ram[60][131]=1;ram[60][132]=0;ram[60][133]=0;ram[60][134]=0;ram[60][135]=0;ram[60][136]=1;
        ram[61][0]=1;ram[61][1]=0;ram[61][2]=1;ram[61][3]=0;ram[61][4]=1;ram[61][5]=0;ram[61][6]=1;ram[61][7]=1;ram[61][8]=0;ram[61][9]=1;ram[61][10]=1;ram[61][11]=0;ram[61][12]=0;ram[61][13]=1;ram[61][14]=1;ram[61][15]=0;ram[61][16]=1;ram[61][17]=0;ram[61][18]=1;ram[61][19]=1;ram[61][20]=1;ram[61][21]=1;ram[61][22]=1;ram[61][23]=1;ram[61][24]=1;ram[61][25]=1;ram[61][26]=1;ram[61][27]=0;ram[61][28]=1;ram[61][29]=1;ram[61][30]=1;ram[61][31]=1;ram[61][32]=1;ram[61][33]=1;ram[61][34]=1;ram[61][35]=0;ram[61][36]=1;ram[61][37]=1;ram[61][38]=1;ram[61][39]=1;ram[61][40]=0;ram[61][41]=0;ram[61][42]=1;ram[61][43]=1;ram[61][44]=0;ram[61][45]=1;ram[61][46]=0;ram[61][47]=1;ram[61][48]=0;ram[61][49]=0;ram[61][50]=1;ram[61][51]=1;ram[61][52]=1;ram[61][53]=0;ram[61][54]=0;ram[61][55]=1;ram[61][56]=1;ram[61][57]=1;ram[61][58]=1;ram[61][59]=1;ram[61][60]=1;ram[61][61]=1;ram[61][62]=1;ram[61][63]=1;ram[61][64]=0;ram[61][65]=1;ram[61][66]=0;ram[61][67]=1;ram[61][68]=1;ram[61][69]=1;ram[61][70]=0;ram[61][71]=1;ram[61][72]=0;ram[61][73]=0;ram[61][74]=1;ram[61][75]=1;ram[61][76]=0;ram[61][77]=1;ram[61][78]=1;ram[61][79]=0;ram[61][80]=1;ram[61][81]=1;ram[61][82]=0;ram[61][83]=1;ram[61][84]=1;ram[61][85]=0;ram[61][86]=1;ram[61][87]=0;ram[61][88]=1;ram[61][89]=0;ram[61][90]=1;ram[61][91]=1;ram[61][92]=1;ram[61][93]=1;ram[61][94]=1;ram[61][95]=0;ram[61][96]=1;ram[61][97]=0;ram[61][98]=1;ram[61][99]=1;ram[61][100]=1;ram[61][101]=1;ram[61][102]=0;ram[61][103]=0;ram[61][104]=1;ram[61][105]=1;ram[61][106]=0;ram[61][107]=1;ram[61][108]=0;ram[61][109]=1;ram[61][110]=1;ram[61][111]=0;ram[61][112]=0;ram[61][113]=1;ram[61][114]=1;ram[61][115]=0;ram[61][116]=1;ram[61][117]=0;ram[61][118]=1;ram[61][119]=0;ram[61][120]=0;ram[61][121]=0;ram[61][122]=0;ram[61][123]=1;ram[61][124]=0;ram[61][125]=0;ram[61][126]=0;ram[61][127]=1;ram[61][128]=1;ram[61][129]=0;ram[61][130]=1;ram[61][131]=1;ram[61][132]=1;ram[61][133]=0;ram[61][134]=1;ram[61][135]=1;ram[61][136]=0;
        ram[62][0]=1;ram[62][1]=1;ram[62][2]=1;ram[62][3]=1;ram[62][4]=0;ram[62][5]=1;ram[62][6]=1;ram[62][7]=1;ram[62][8]=0;ram[62][9]=0;ram[62][10]=1;ram[62][11]=0;ram[62][12]=1;ram[62][13]=0;ram[62][14]=1;ram[62][15]=1;ram[62][16]=1;ram[62][17]=0;ram[62][18]=1;ram[62][19]=0;ram[62][20]=1;ram[62][21]=1;ram[62][22]=1;ram[62][23]=1;ram[62][24]=1;ram[62][25]=1;ram[62][26]=1;ram[62][27]=1;ram[62][28]=1;ram[62][29]=1;ram[62][30]=1;ram[62][31]=1;ram[62][32]=1;ram[62][33]=1;ram[62][34]=1;ram[62][35]=0;ram[62][36]=1;ram[62][37]=1;ram[62][38]=0;ram[62][39]=1;ram[62][40]=1;ram[62][41]=1;ram[62][42]=0;ram[62][43]=1;ram[62][44]=1;ram[62][45]=0;ram[62][46]=1;ram[62][47]=1;ram[62][48]=1;ram[62][49]=1;ram[62][50]=1;ram[62][51]=1;ram[62][52]=1;ram[62][53]=0;ram[62][54]=0;ram[62][55]=0;ram[62][56]=0;ram[62][57]=0;ram[62][58]=1;ram[62][59]=1;ram[62][60]=0;ram[62][61]=1;ram[62][62]=1;ram[62][63]=1;ram[62][64]=1;ram[62][65]=1;ram[62][66]=1;ram[62][67]=1;ram[62][68]=1;ram[62][69]=0;ram[62][70]=0;ram[62][71]=1;ram[62][72]=1;ram[62][73]=1;ram[62][74]=0;ram[62][75]=1;ram[62][76]=0;ram[62][77]=1;ram[62][78]=0;ram[62][79]=1;ram[62][80]=1;ram[62][81]=1;ram[62][82]=1;ram[62][83]=0;ram[62][84]=1;ram[62][85]=1;ram[62][86]=0;ram[62][87]=1;ram[62][88]=1;ram[62][89]=1;ram[62][90]=1;ram[62][91]=1;ram[62][92]=0;ram[62][93]=1;ram[62][94]=1;ram[62][95]=0;ram[62][96]=1;ram[62][97]=0;ram[62][98]=1;ram[62][99]=0;ram[62][100]=0;ram[62][101]=1;ram[62][102]=1;ram[62][103]=1;ram[62][104]=1;ram[62][105]=0;ram[62][106]=1;ram[62][107]=1;ram[62][108]=0;ram[62][109]=1;ram[62][110]=1;ram[62][111]=0;ram[62][112]=1;ram[62][113]=1;ram[62][114]=1;ram[62][115]=1;ram[62][116]=1;ram[62][117]=1;ram[62][118]=1;ram[62][119]=1;ram[62][120]=1;ram[62][121]=0;ram[62][122]=1;ram[62][123]=1;ram[62][124]=0;ram[62][125]=0;ram[62][126]=1;ram[62][127]=0;ram[62][128]=1;ram[62][129]=1;ram[62][130]=1;ram[62][131]=0;ram[62][132]=0;ram[62][133]=0;ram[62][134]=1;ram[62][135]=1;ram[62][136]=1;
        ram[63][0]=1;ram[63][1]=1;ram[63][2]=0;ram[63][3]=1;ram[63][4]=0;ram[63][5]=0;ram[63][6]=1;ram[63][7]=1;ram[63][8]=1;ram[63][9]=1;ram[63][10]=0;ram[63][11]=0;ram[63][12]=0;ram[63][13]=1;ram[63][14]=0;ram[63][15]=1;ram[63][16]=0;ram[63][17]=1;ram[63][18]=0;ram[63][19]=0;ram[63][20]=1;ram[63][21]=1;ram[63][22]=1;ram[63][23]=1;ram[63][24]=1;ram[63][25]=1;ram[63][26]=0;ram[63][27]=0;ram[63][28]=1;ram[63][29]=1;ram[63][30]=1;ram[63][31]=1;ram[63][32]=0;ram[63][33]=0;ram[63][34]=1;ram[63][35]=0;ram[63][36]=1;ram[63][37]=1;ram[63][38]=0;ram[63][39]=1;ram[63][40]=0;ram[63][41]=0;ram[63][42]=1;ram[63][43]=1;ram[63][44]=1;ram[63][45]=0;ram[63][46]=0;ram[63][47]=1;ram[63][48]=1;ram[63][49]=1;ram[63][50]=1;ram[63][51]=1;ram[63][52]=0;ram[63][53]=0;ram[63][54]=1;ram[63][55]=0;ram[63][56]=1;ram[63][57]=0;ram[63][58]=0;ram[63][59]=1;ram[63][60]=1;ram[63][61]=1;ram[63][62]=1;ram[63][63]=0;ram[63][64]=1;ram[63][65]=1;ram[63][66]=1;ram[63][67]=0;ram[63][68]=0;ram[63][69]=1;ram[63][70]=0;ram[63][71]=0;ram[63][72]=1;ram[63][73]=0;ram[63][74]=0;ram[63][75]=1;ram[63][76]=0;ram[63][77]=1;ram[63][78]=1;ram[63][79]=1;ram[63][80]=1;ram[63][81]=0;ram[63][82]=0;ram[63][83]=1;ram[63][84]=1;ram[63][85]=0;ram[63][86]=1;ram[63][87]=1;ram[63][88]=1;ram[63][89]=1;ram[63][90]=0;ram[63][91]=1;ram[63][92]=0;ram[63][93]=1;ram[63][94]=1;ram[63][95]=1;ram[63][96]=1;ram[63][97]=0;ram[63][98]=0;ram[63][99]=1;ram[63][100]=0;ram[63][101]=0;ram[63][102]=1;ram[63][103]=1;ram[63][104]=0;ram[63][105]=1;ram[63][106]=1;ram[63][107]=1;ram[63][108]=1;ram[63][109]=0;ram[63][110]=1;ram[63][111]=1;ram[63][112]=0;ram[63][113]=0;ram[63][114]=1;ram[63][115]=1;ram[63][116]=0;ram[63][117]=0;ram[63][118]=1;ram[63][119]=1;ram[63][120]=0;ram[63][121]=0;ram[63][122]=0;ram[63][123]=0;ram[63][124]=0;ram[63][125]=1;ram[63][126]=1;ram[63][127]=1;ram[63][128]=1;ram[63][129]=1;ram[63][130]=0;ram[63][131]=0;ram[63][132]=0;ram[63][133]=0;ram[63][134]=1;ram[63][135]=1;ram[63][136]=0;
        ram[64][0]=1;ram[64][1]=1;ram[64][2]=1;ram[64][3]=1;ram[64][4]=1;ram[64][5]=1;ram[64][6]=1;ram[64][7]=1;ram[64][8]=0;ram[64][9]=0;ram[64][10]=0;ram[64][11]=0;ram[64][12]=0;ram[64][13]=1;ram[64][14]=1;ram[64][15]=0;ram[64][16]=1;ram[64][17]=0;ram[64][18]=1;ram[64][19]=0;ram[64][20]=1;ram[64][21]=1;ram[64][22]=0;ram[64][23]=0;ram[64][24]=1;ram[64][25]=1;ram[64][26]=1;ram[64][27]=0;ram[64][28]=0;ram[64][29]=0;ram[64][30]=0;ram[64][31]=0;ram[64][32]=1;ram[64][33]=1;ram[64][34]=1;ram[64][35]=1;ram[64][36]=1;ram[64][37]=1;ram[64][38]=1;ram[64][39]=1;ram[64][40]=0;ram[64][41]=1;ram[64][42]=1;ram[64][43]=1;ram[64][44]=0;ram[64][45]=1;ram[64][46]=1;ram[64][47]=1;ram[64][48]=1;ram[64][49]=0;ram[64][50]=1;ram[64][51]=1;ram[64][52]=1;ram[64][53]=1;ram[64][54]=0;ram[64][55]=1;ram[64][56]=1;ram[64][57]=0;ram[64][58]=1;ram[64][59]=1;ram[64][60]=0;ram[64][61]=1;ram[64][62]=1;ram[64][63]=1;ram[64][64]=0;ram[64][65]=0;ram[64][66]=1;ram[64][67]=1;ram[64][68]=1;ram[64][69]=0;ram[64][70]=0;ram[64][71]=0;ram[64][72]=1;ram[64][73]=1;ram[64][74]=0;ram[64][75]=1;ram[64][76]=0;ram[64][77]=1;ram[64][78]=0;ram[64][79]=1;ram[64][80]=1;ram[64][81]=1;ram[64][82]=0;ram[64][83]=1;ram[64][84]=1;ram[64][85]=1;ram[64][86]=0;ram[64][87]=1;ram[64][88]=0;ram[64][89]=0;ram[64][90]=1;ram[64][91]=0;ram[64][92]=1;ram[64][93]=0;ram[64][94]=1;ram[64][95]=1;ram[64][96]=1;ram[64][97]=0;ram[64][98]=0;ram[64][99]=1;ram[64][100]=1;ram[64][101]=0;ram[64][102]=0;ram[64][103]=1;ram[64][104]=1;ram[64][105]=1;ram[64][106]=0;ram[64][107]=1;ram[64][108]=0;ram[64][109]=1;ram[64][110]=1;ram[64][111]=1;ram[64][112]=1;ram[64][113]=0;ram[64][114]=0;ram[64][115]=0;ram[64][116]=1;ram[64][117]=1;ram[64][118]=0;ram[64][119]=0;ram[64][120]=0;ram[64][121]=0;ram[64][122]=1;ram[64][123]=1;ram[64][124]=1;ram[64][125]=1;ram[64][126]=1;ram[64][127]=1;ram[64][128]=0;ram[64][129]=0;ram[64][130]=1;ram[64][131]=1;ram[64][132]=0;ram[64][133]=0;ram[64][134]=1;ram[64][135]=1;ram[64][136]=0;
        ram[65][0]=0;ram[65][1]=1;ram[65][2]=0;ram[65][3]=1;ram[65][4]=1;ram[65][5]=0;ram[65][6]=1;ram[65][7]=1;ram[65][8]=1;ram[65][9]=0;ram[65][10]=0;ram[65][11]=1;ram[65][12]=1;ram[65][13]=1;ram[65][14]=0;ram[65][15]=0;ram[65][16]=1;ram[65][17]=0;ram[65][18]=1;ram[65][19]=0;ram[65][20]=0;ram[65][21]=0;ram[65][22]=1;ram[65][23]=1;ram[65][24]=1;ram[65][25]=1;ram[65][26]=1;ram[65][27]=1;ram[65][28]=0;ram[65][29]=1;ram[65][30]=0;ram[65][31]=0;ram[65][32]=0;ram[65][33]=1;ram[65][34]=1;ram[65][35]=1;ram[65][36]=1;ram[65][37]=0;ram[65][38]=1;ram[65][39]=1;ram[65][40]=1;ram[65][41]=1;ram[65][42]=1;ram[65][43]=1;ram[65][44]=0;ram[65][45]=0;ram[65][46]=1;ram[65][47]=1;ram[65][48]=1;ram[65][49]=0;ram[65][50]=1;ram[65][51]=0;ram[65][52]=1;ram[65][53]=1;ram[65][54]=0;ram[65][55]=1;ram[65][56]=0;ram[65][57]=0;ram[65][58]=0;ram[65][59]=1;ram[65][60]=1;ram[65][61]=0;ram[65][62]=0;ram[65][63]=1;ram[65][64]=1;ram[65][65]=1;ram[65][66]=0;ram[65][67]=1;ram[65][68]=1;ram[65][69]=0;ram[65][70]=1;ram[65][71]=1;ram[65][72]=1;ram[65][73]=0;ram[65][74]=0;ram[65][75]=0;ram[65][76]=1;ram[65][77]=0;ram[65][78]=0;ram[65][79]=1;ram[65][80]=1;ram[65][81]=0;ram[65][82]=1;ram[65][83]=1;ram[65][84]=1;ram[65][85]=0;ram[65][86]=0;ram[65][87]=1;ram[65][88]=1;ram[65][89]=1;ram[65][90]=0;ram[65][91]=1;ram[65][92]=0;ram[65][93]=1;ram[65][94]=1;ram[65][95]=0;ram[65][96]=1;ram[65][97]=1;ram[65][98]=1;ram[65][99]=1;ram[65][100]=1;ram[65][101]=0;ram[65][102]=1;ram[65][103]=1;ram[65][104]=1;ram[65][105]=1;ram[65][106]=1;ram[65][107]=0;ram[65][108]=0;ram[65][109]=1;ram[65][110]=0;ram[65][111]=1;ram[65][112]=0;ram[65][113]=1;ram[65][114]=0;ram[65][115]=1;ram[65][116]=1;ram[65][117]=0;ram[65][118]=0;ram[65][119]=0;ram[65][120]=0;ram[65][121]=0;ram[65][122]=0;ram[65][123]=1;ram[65][124]=0;ram[65][125]=1;ram[65][126]=0;ram[65][127]=1;ram[65][128]=0;ram[65][129]=1;ram[65][130]=1;ram[65][131]=0;ram[65][132]=0;ram[65][133]=1;ram[65][134]=1;ram[65][135]=1;ram[65][136]=1;
        ram[66][0]=1;ram[66][1]=1;ram[66][2]=1;ram[66][3]=1;ram[66][4]=1;ram[66][5]=1;ram[66][6]=0;ram[66][7]=1;ram[66][8]=1;ram[66][9]=1;ram[66][10]=0;ram[66][11]=1;ram[66][12]=0;ram[66][13]=0;ram[66][14]=1;ram[66][15]=1;ram[66][16]=1;ram[66][17]=1;ram[66][18]=1;ram[66][19]=1;ram[66][20]=0;ram[66][21]=1;ram[66][22]=1;ram[66][23]=1;ram[66][24]=1;ram[66][25]=0;ram[66][26]=1;ram[66][27]=1;ram[66][28]=1;ram[66][29]=1;ram[66][30]=1;ram[66][31]=0;ram[66][32]=1;ram[66][33]=0;ram[66][34]=1;ram[66][35]=0;ram[66][36]=1;ram[66][37]=0;ram[66][38]=0;ram[66][39]=1;ram[66][40]=1;ram[66][41]=0;ram[66][42]=1;ram[66][43]=0;ram[66][44]=0;ram[66][45]=0;ram[66][46]=1;ram[66][47]=0;ram[66][48]=1;ram[66][49]=1;ram[66][50]=1;ram[66][51]=1;ram[66][52]=1;ram[66][53]=1;ram[66][54]=1;ram[66][55]=1;ram[66][56]=1;ram[66][57]=1;ram[66][58]=0;ram[66][59]=1;ram[66][60]=1;ram[66][61]=1;ram[66][62]=1;ram[66][63]=0;ram[66][64]=0;ram[66][65]=0;ram[66][66]=0;ram[66][67]=1;ram[66][68]=1;ram[66][69]=1;ram[66][70]=1;ram[66][71]=1;ram[66][72]=1;ram[66][73]=1;ram[66][74]=1;ram[66][75]=1;ram[66][76]=0;ram[66][77]=1;ram[66][78]=1;ram[66][79]=0;ram[66][80]=1;ram[66][81]=1;ram[66][82]=0;ram[66][83]=0;ram[66][84]=0;ram[66][85]=0;ram[66][86]=1;ram[66][87]=0;ram[66][88]=1;ram[66][89]=0;ram[66][90]=1;ram[66][91]=1;ram[66][92]=0;ram[66][93]=1;ram[66][94]=1;ram[66][95]=1;ram[66][96]=1;ram[66][97]=0;ram[66][98]=1;ram[66][99]=0;ram[66][100]=1;ram[66][101]=0;ram[66][102]=1;ram[66][103]=1;ram[66][104]=0;ram[66][105]=1;ram[66][106]=1;ram[66][107]=1;ram[66][108]=1;ram[66][109]=1;ram[66][110]=0;ram[66][111]=0;ram[66][112]=0;ram[66][113]=0;ram[66][114]=1;ram[66][115]=0;ram[66][116]=0;ram[66][117]=1;ram[66][118]=0;ram[66][119]=0;ram[66][120]=1;ram[66][121]=1;ram[66][122]=1;ram[66][123]=1;ram[66][124]=1;ram[66][125]=0;ram[66][126]=1;ram[66][127]=1;ram[66][128]=1;ram[66][129]=1;ram[66][130]=1;ram[66][131]=1;ram[66][132]=1;ram[66][133]=0;ram[66][134]=1;ram[66][135]=1;ram[66][136]=0;
        ram[67][0]=1;ram[67][1]=1;ram[67][2]=0;ram[67][3]=1;ram[67][4]=1;ram[67][5]=1;ram[67][6]=0;ram[67][7]=0;ram[67][8]=1;ram[67][9]=1;ram[67][10]=0;ram[67][11]=1;ram[67][12]=1;ram[67][13]=0;ram[67][14]=1;ram[67][15]=1;ram[67][16]=1;ram[67][17]=0;ram[67][18]=0;ram[67][19]=0;ram[67][20]=1;ram[67][21]=0;ram[67][22]=0;ram[67][23]=0;ram[67][24]=0;ram[67][25]=0;ram[67][26]=1;ram[67][27]=1;ram[67][28]=1;ram[67][29]=1;ram[67][30]=1;ram[67][31]=1;ram[67][32]=1;ram[67][33]=1;ram[67][34]=1;ram[67][35]=0;ram[67][36]=1;ram[67][37]=1;ram[67][38]=0;ram[67][39]=1;ram[67][40]=1;ram[67][41]=0;ram[67][42]=1;ram[67][43]=0;ram[67][44]=1;ram[67][45]=1;ram[67][46]=1;ram[67][47]=1;ram[67][48]=1;ram[67][49]=1;ram[67][50]=1;ram[67][51]=1;ram[67][52]=1;ram[67][53]=0;ram[67][54]=1;ram[67][55]=0;ram[67][56]=1;ram[67][57]=1;ram[67][58]=0;ram[67][59]=1;ram[67][60]=1;ram[67][61]=0;ram[67][62]=0;ram[67][63]=1;ram[67][64]=0;ram[67][65]=0;ram[67][66]=0;ram[67][67]=1;ram[67][68]=1;ram[67][69]=0;ram[67][70]=1;ram[67][71]=0;ram[67][72]=1;ram[67][73]=1;ram[67][74]=1;ram[67][75]=1;ram[67][76]=1;ram[67][77]=1;ram[67][78]=1;ram[67][79]=0;ram[67][80]=1;ram[67][81]=1;ram[67][82]=1;ram[67][83]=1;ram[67][84]=1;ram[67][85]=0;ram[67][86]=1;ram[67][87]=1;ram[67][88]=1;ram[67][89]=0;ram[67][90]=0;ram[67][91]=0;ram[67][92]=1;ram[67][93]=1;ram[67][94]=0;ram[67][95]=1;ram[67][96]=1;ram[67][97]=0;ram[67][98]=1;ram[67][99]=1;ram[67][100]=1;ram[67][101]=1;ram[67][102]=1;ram[67][103]=1;ram[67][104]=1;ram[67][105]=0;ram[67][106]=1;ram[67][107]=1;ram[67][108]=0;ram[67][109]=1;ram[67][110]=0;ram[67][111]=1;ram[67][112]=0;ram[67][113]=1;ram[67][114]=1;ram[67][115]=1;ram[67][116]=1;ram[67][117]=1;ram[67][118]=0;ram[67][119]=1;ram[67][120]=1;ram[67][121]=0;ram[67][122]=0;ram[67][123]=1;ram[67][124]=1;ram[67][125]=1;ram[67][126]=1;ram[67][127]=0;ram[67][128]=1;ram[67][129]=0;ram[67][130]=1;ram[67][131]=0;ram[67][132]=1;ram[67][133]=1;ram[67][134]=1;ram[67][135]=0;ram[67][136]=1;
        ram[68][0]=1;ram[68][1]=1;ram[68][2]=1;ram[68][3]=1;ram[68][4]=1;ram[68][5]=1;ram[68][6]=1;ram[68][7]=0;ram[68][8]=1;ram[68][9]=0;ram[68][10]=1;ram[68][11]=1;ram[68][12]=1;ram[68][13]=0;ram[68][14]=1;ram[68][15]=0;ram[68][16]=1;ram[68][17]=0;ram[68][18]=1;ram[68][19]=1;ram[68][20]=1;ram[68][21]=1;ram[68][22]=0;ram[68][23]=1;ram[68][24]=0;ram[68][25]=0;ram[68][26]=1;ram[68][27]=1;ram[68][28]=1;ram[68][29]=0;ram[68][30]=0;ram[68][31]=0;ram[68][32]=0;ram[68][33]=1;ram[68][34]=0;ram[68][35]=0;ram[68][36]=0;ram[68][37]=0;ram[68][38]=0;ram[68][39]=0;ram[68][40]=0;ram[68][41]=0;ram[68][42]=0;ram[68][43]=0;ram[68][44]=1;ram[68][45]=0;ram[68][46]=1;ram[68][47]=0;ram[68][48]=0;ram[68][49]=1;ram[68][50]=1;ram[68][51]=0;ram[68][52]=1;ram[68][53]=0;ram[68][54]=1;ram[68][55]=1;ram[68][56]=1;ram[68][57]=1;ram[68][58]=0;ram[68][59]=1;ram[68][60]=0;ram[68][61]=1;ram[68][62]=1;ram[68][63]=1;ram[68][64]=0;ram[68][65]=0;ram[68][66]=0;ram[68][67]=1;ram[68][68]=0;ram[68][69]=0;ram[68][70]=0;ram[68][71]=1;ram[68][72]=0;ram[68][73]=0;ram[68][74]=0;ram[68][75]=0;ram[68][76]=1;ram[68][77]=0;ram[68][78]=0;ram[68][79]=1;ram[68][80]=0;ram[68][81]=0;ram[68][82]=1;ram[68][83]=0;ram[68][84]=0;ram[68][85]=1;ram[68][86]=1;ram[68][87]=0;ram[68][88]=1;ram[68][89]=1;ram[68][90]=1;ram[68][91]=0;ram[68][92]=1;ram[68][93]=1;ram[68][94]=0;ram[68][95]=1;ram[68][96]=1;ram[68][97]=0;ram[68][98]=1;ram[68][99]=0;ram[68][100]=0;ram[68][101]=0;ram[68][102]=1;ram[68][103]=1;ram[68][104]=1;ram[68][105]=0;ram[68][106]=1;ram[68][107]=0;ram[68][108]=1;ram[68][109]=1;ram[68][110]=1;ram[68][111]=1;ram[68][112]=1;ram[68][113]=0;ram[68][114]=1;ram[68][115]=1;ram[68][116]=1;ram[68][117]=0;ram[68][118]=1;ram[68][119]=1;ram[68][120]=0;ram[68][121]=1;ram[68][122]=0;ram[68][123]=1;ram[68][124]=0;ram[68][125]=0;ram[68][126]=0;ram[68][127]=0;ram[68][128]=1;ram[68][129]=1;ram[68][130]=1;ram[68][131]=1;ram[68][132]=1;ram[68][133]=0;ram[68][134]=1;ram[68][135]=1;ram[68][136]=1;
        ram[69][0]=1;ram[69][1]=1;ram[69][2]=1;ram[69][3]=1;ram[69][4]=0;ram[69][5]=0;ram[69][6]=1;ram[69][7]=1;ram[69][8]=1;ram[69][9]=1;ram[69][10]=1;ram[69][11]=0;ram[69][12]=1;ram[69][13]=0;ram[69][14]=0;ram[69][15]=1;ram[69][16]=1;ram[69][17]=1;ram[69][18]=1;ram[69][19]=0;ram[69][20]=1;ram[69][21]=0;ram[69][22]=1;ram[69][23]=0;ram[69][24]=0;ram[69][25]=1;ram[69][26]=0;ram[69][27]=0;ram[69][28]=1;ram[69][29]=1;ram[69][30]=1;ram[69][31]=1;ram[69][32]=1;ram[69][33]=1;ram[69][34]=0;ram[69][35]=1;ram[69][36]=0;ram[69][37]=1;ram[69][38]=1;ram[69][39]=1;ram[69][40]=1;ram[69][41]=1;ram[69][42]=1;ram[69][43]=1;ram[69][44]=1;ram[69][45]=1;ram[69][46]=0;ram[69][47]=1;ram[69][48]=1;ram[69][49]=1;ram[69][50]=1;ram[69][51]=1;ram[69][52]=0;ram[69][53]=1;ram[69][54]=1;ram[69][55]=0;ram[69][56]=0;ram[69][57]=1;ram[69][58]=1;ram[69][59]=1;ram[69][60]=1;ram[69][61]=0;ram[69][62]=1;ram[69][63]=1;ram[69][64]=0;ram[69][65]=0;ram[69][66]=1;ram[69][67]=1;ram[69][68]=1;ram[69][69]=1;ram[69][70]=1;ram[69][71]=1;ram[69][72]=0;ram[69][73]=1;ram[69][74]=1;ram[69][75]=1;ram[69][76]=0;ram[69][77]=0;ram[69][78]=0;ram[69][79]=1;ram[69][80]=1;ram[69][81]=1;ram[69][82]=1;ram[69][83]=1;ram[69][84]=1;ram[69][85]=0;ram[69][86]=1;ram[69][87]=0;ram[69][88]=1;ram[69][89]=0;ram[69][90]=1;ram[69][91]=1;ram[69][92]=1;ram[69][93]=1;ram[69][94]=1;ram[69][95]=0;ram[69][96]=1;ram[69][97]=1;ram[69][98]=1;ram[69][99]=1;ram[69][100]=1;ram[69][101]=1;ram[69][102]=1;ram[69][103]=1;ram[69][104]=1;ram[69][105]=1;ram[69][106]=1;ram[69][107]=0;ram[69][108]=0;ram[69][109]=1;ram[69][110]=1;ram[69][111]=0;ram[69][112]=0;ram[69][113]=1;ram[69][114]=0;ram[69][115]=0;ram[69][116]=1;ram[69][117]=1;ram[69][118]=0;ram[69][119]=0;ram[69][120]=0;ram[69][121]=1;ram[69][122]=1;ram[69][123]=0;ram[69][124]=0;ram[69][125]=0;ram[69][126]=0;ram[69][127]=1;ram[69][128]=1;ram[69][129]=0;ram[69][130]=1;ram[69][131]=0;ram[69][132]=1;ram[69][133]=1;ram[69][134]=1;ram[69][135]=0;ram[69][136]=0;
        ram[70][0]=1;ram[70][1]=1;ram[70][2]=0;ram[70][3]=1;ram[70][4]=1;ram[70][5]=1;ram[70][6]=0;ram[70][7]=0;ram[70][8]=0;ram[70][9]=0;ram[70][10]=1;ram[70][11]=0;ram[70][12]=1;ram[70][13]=1;ram[70][14]=0;ram[70][15]=1;ram[70][16]=1;ram[70][17]=0;ram[70][18]=1;ram[70][19]=1;ram[70][20]=0;ram[70][21]=0;ram[70][22]=1;ram[70][23]=0;ram[70][24]=0;ram[70][25]=0;ram[70][26]=0;ram[70][27]=0;ram[70][28]=0;ram[70][29]=1;ram[70][30]=0;ram[70][31]=1;ram[70][32]=1;ram[70][33]=1;ram[70][34]=1;ram[70][35]=1;ram[70][36]=1;ram[70][37]=1;ram[70][38]=0;ram[70][39]=0;ram[70][40]=1;ram[70][41]=1;ram[70][42]=1;ram[70][43]=1;ram[70][44]=1;ram[70][45]=1;ram[70][46]=1;ram[70][47]=1;ram[70][48]=1;ram[70][49]=1;ram[70][50]=1;ram[70][51]=1;ram[70][52]=0;ram[70][53]=1;ram[70][54]=0;ram[70][55]=0;ram[70][56]=1;ram[70][57]=1;ram[70][58]=1;ram[70][59]=1;ram[70][60]=1;ram[70][61]=1;ram[70][62]=1;ram[70][63]=0;ram[70][64]=0;ram[70][65]=1;ram[70][66]=1;ram[70][67]=1;ram[70][68]=1;ram[70][69]=1;ram[70][70]=0;ram[70][71]=0;ram[70][72]=1;ram[70][73]=1;ram[70][74]=1;ram[70][75]=1;ram[70][76]=0;ram[70][77]=1;ram[70][78]=1;ram[70][79]=1;ram[70][80]=0;ram[70][81]=0;ram[70][82]=1;ram[70][83]=1;ram[70][84]=1;ram[70][85]=1;ram[70][86]=1;ram[70][87]=0;ram[70][88]=1;ram[70][89]=0;ram[70][90]=0;ram[70][91]=1;ram[70][92]=1;ram[70][93]=0;ram[70][94]=1;ram[70][95]=1;ram[70][96]=1;ram[70][97]=1;ram[70][98]=1;ram[70][99]=1;ram[70][100]=1;ram[70][101]=1;ram[70][102]=1;ram[70][103]=1;ram[70][104]=1;ram[70][105]=0;ram[70][106]=1;ram[70][107]=0;ram[70][108]=1;ram[70][109]=1;ram[70][110]=1;ram[70][111]=1;ram[70][112]=1;ram[70][113]=0;ram[70][114]=1;ram[70][115]=1;ram[70][116]=1;ram[70][117]=0;ram[70][118]=1;ram[70][119]=0;ram[70][120]=1;ram[70][121]=0;ram[70][122]=0;ram[70][123]=1;ram[70][124]=0;ram[70][125]=1;ram[70][126]=1;ram[70][127]=1;ram[70][128]=0;ram[70][129]=0;ram[70][130]=1;ram[70][131]=1;ram[70][132]=0;ram[70][133]=1;ram[70][134]=1;ram[70][135]=0;ram[70][136]=1;
        ram[71][0]=1;ram[71][1]=1;ram[71][2]=1;ram[71][3]=0;ram[71][4]=0;ram[71][5]=1;ram[71][6]=1;ram[71][7]=0;ram[71][8]=1;ram[71][9]=0;ram[71][10]=1;ram[71][11]=1;ram[71][12]=0;ram[71][13]=0;ram[71][14]=1;ram[71][15]=1;ram[71][16]=0;ram[71][17]=0;ram[71][18]=1;ram[71][19]=0;ram[71][20]=0;ram[71][21]=1;ram[71][22]=1;ram[71][23]=1;ram[71][24]=1;ram[71][25]=1;ram[71][26]=1;ram[71][27]=0;ram[71][28]=0;ram[71][29]=1;ram[71][30]=0;ram[71][31]=0;ram[71][32]=1;ram[71][33]=1;ram[71][34]=0;ram[71][35]=1;ram[71][36]=1;ram[71][37]=1;ram[71][38]=1;ram[71][39]=1;ram[71][40]=0;ram[71][41]=1;ram[71][42]=0;ram[71][43]=0;ram[71][44]=1;ram[71][45]=0;ram[71][46]=1;ram[71][47]=1;ram[71][48]=1;ram[71][49]=1;ram[71][50]=1;ram[71][51]=1;ram[71][52]=1;ram[71][53]=1;ram[71][54]=0;ram[71][55]=1;ram[71][56]=1;ram[71][57]=1;ram[71][58]=1;ram[71][59]=0;ram[71][60]=0;ram[71][61]=1;ram[71][62]=1;ram[71][63]=1;ram[71][64]=0;ram[71][65]=0;ram[71][66]=0;ram[71][67]=0;ram[71][68]=0;ram[71][69]=1;ram[71][70]=0;ram[71][71]=1;ram[71][72]=1;ram[71][73]=1;ram[71][74]=1;ram[71][75]=0;ram[71][76]=1;ram[71][77]=1;ram[71][78]=0;ram[71][79]=1;ram[71][80]=0;ram[71][81]=1;ram[71][82]=0;ram[71][83]=1;ram[71][84]=0;ram[71][85]=0;ram[71][86]=0;ram[71][87]=0;ram[71][88]=1;ram[71][89]=1;ram[71][90]=1;ram[71][91]=0;ram[71][92]=0;ram[71][93]=1;ram[71][94]=0;ram[71][95]=1;ram[71][96]=1;ram[71][97]=1;ram[71][98]=0;ram[71][99]=0;ram[71][100]=0;ram[71][101]=1;ram[71][102]=0;ram[71][103]=1;ram[71][104]=1;ram[71][105]=1;ram[71][106]=1;ram[71][107]=1;ram[71][108]=1;ram[71][109]=1;ram[71][110]=1;ram[71][111]=0;ram[71][112]=1;ram[71][113]=1;ram[71][114]=0;ram[71][115]=0;ram[71][116]=0;ram[71][117]=1;ram[71][118]=0;ram[71][119]=1;ram[71][120]=1;ram[71][121]=0;ram[71][122]=0;ram[71][123]=1;ram[71][124]=1;ram[71][125]=0;ram[71][126]=1;ram[71][127]=1;ram[71][128]=1;ram[71][129]=1;ram[71][130]=1;ram[71][131]=1;ram[71][132]=0;ram[71][133]=1;ram[71][134]=1;ram[71][135]=1;ram[71][136]=0;
        ram[72][0]=1;ram[72][1]=0;ram[72][2]=0;ram[72][3]=1;ram[72][4]=1;ram[72][5]=1;ram[72][6]=1;ram[72][7]=1;ram[72][8]=0;ram[72][9]=0;ram[72][10]=1;ram[72][11]=0;ram[72][12]=1;ram[72][13]=0;ram[72][14]=0;ram[72][15]=1;ram[72][16]=1;ram[72][17]=1;ram[72][18]=1;ram[72][19]=1;ram[72][20]=1;ram[72][21]=0;ram[72][22]=0;ram[72][23]=1;ram[72][24]=1;ram[72][25]=1;ram[72][26]=1;ram[72][27]=0;ram[72][28]=1;ram[72][29]=1;ram[72][30]=1;ram[72][31]=1;ram[72][32]=1;ram[72][33]=1;ram[72][34]=1;ram[72][35]=1;ram[72][36]=1;ram[72][37]=1;ram[72][38]=1;ram[72][39]=1;ram[72][40]=1;ram[72][41]=0;ram[72][42]=0;ram[72][43]=1;ram[72][44]=0;ram[72][45]=1;ram[72][46]=1;ram[72][47]=1;ram[72][48]=1;ram[72][49]=0;ram[72][50]=0;ram[72][51]=0;ram[72][52]=1;ram[72][53]=1;ram[72][54]=1;ram[72][55]=1;ram[72][56]=1;ram[72][57]=1;ram[72][58]=1;ram[72][59]=0;ram[72][60]=1;ram[72][61]=0;ram[72][62]=1;ram[72][63]=1;ram[72][64]=1;ram[72][65]=1;ram[72][66]=1;ram[72][67]=1;ram[72][68]=1;ram[72][69]=0;ram[72][70]=1;ram[72][71]=0;ram[72][72]=1;ram[72][73]=1;ram[72][74]=0;ram[72][75]=1;ram[72][76]=1;ram[72][77]=0;ram[72][78]=1;ram[72][79]=0;ram[72][80]=0;ram[72][81]=1;ram[72][82]=0;ram[72][83]=0;ram[72][84]=1;ram[72][85]=1;ram[72][86]=1;ram[72][87]=1;ram[72][88]=1;ram[72][89]=1;ram[72][90]=0;ram[72][91]=0;ram[72][92]=0;ram[72][93]=1;ram[72][94]=1;ram[72][95]=1;ram[72][96]=0;ram[72][97]=1;ram[72][98]=1;ram[72][99]=1;ram[72][100]=0;ram[72][101]=1;ram[72][102]=1;ram[72][103]=1;ram[72][104]=1;ram[72][105]=0;ram[72][106]=1;ram[72][107]=1;ram[72][108]=1;ram[72][109]=1;ram[72][110]=1;ram[72][111]=0;ram[72][112]=0;ram[72][113]=1;ram[72][114]=1;ram[72][115]=1;ram[72][116]=0;ram[72][117]=1;ram[72][118]=0;ram[72][119]=1;ram[72][120]=0;ram[72][121]=0;ram[72][122]=0;ram[72][123]=1;ram[72][124]=1;ram[72][125]=1;ram[72][126]=1;ram[72][127]=0;ram[72][128]=0;ram[72][129]=1;ram[72][130]=0;ram[72][131]=1;ram[72][132]=1;ram[72][133]=0;ram[72][134]=1;ram[72][135]=0;ram[72][136]=1;
        ram[73][0]=1;ram[73][1]=1;ram[73][2]=0;ram[73][3]=0;ram[73][4]=1;ram[73][5]=0;ram[73][6]=0;ram[73][7]=1;ram[73][8]=0;ram[73][9]=0;ram[73][10]=1;ram[73][11]=1;ram[73][12]=1;ram[73][13]=1;ram[73][14]=0;ram[73][15]=1;ram[73][16]=0;ram[73][17]=1;ram[73][18]=0;ram[73][19]=1;ram[73][20]=1;ram[73][21]=1;ram[73][22]=1;ram[73][23]=1;ram[73][24]=1;ram[73][25]=1;ram[73][26]=1;ram[73][27]=1;ram[73][28]=0;ram[73][29]=1;ram[73][30]=1;ram[73][31]=1;ram[73][32]=1;ram[73][33]=1;ram[73][34]=0;ram[73][35]=1;ram[73][36]=0;ram[73][37]=1;ram[73][38]=1;ram[73][39]=1;ram[73][40]=0;ram[73][41]=1;ram[73][42]=1;ram[73][43]=0;ram[73][44]=1;ram[73][45]=1;ram[73][46]=0;ram[73][47]=1;ram[73][48]=1;ram[73][49]=0;ram[73][50]=0;ram[73][51]=1;ram[73][52]=0;ram[73][53]=1;ram[73][54]=0;ram[73][55]=0;ram[73][56]=1;ram[73][57]=0;ram[73][58]=1;ram[73][59]=1;ram[73][60]=1;ram[73][61]=1;ram[73][62]=1;ram[73][63]=1;ram[73][64]=1;ram[73][65]=0;ram[73][66]=1;ram[73][67]=0;ram[73][68]=0;ram[73][69]=1;ram[73][70]=0;ram[73][71]=1;ram[73][72]=1;ram[73][73]=0;ram[73][74]=1;ram[73][75]=1;ram[73][76]=1;ram[73][77]=0;ram[73][78]=1;ram[73][79]=0;ram[73][80]=0;ram[73][81]=0;ram[73][82]=1;ram[73][83]=0;ram[73][84]=1;ram[73][85]=0;ram[73][86]=1;ram[73][87]=1;ram[73][88]=1;ram[73][89]=1;ram[73][90]=0;ram[73][91]=1;ram[73][92]=0;ram[73][93]=1;ram[73][94]=1;ram[73][95]=1;ram[73][96]=0;ram[73][97]=1;ram[73][98]=1;ram[73][99]=1;ram[73][100]=1;ram[73][101]=1;ram[73][102]=1;ram[73][103]=1;ram[73][104]=1;ram[73][105]=1;ram[73][106]=1;ram[73][107]=0;ram[73][108]=0;ram[73][109]=0;ram[73][110]=0;ram[73][111]=0;ram[73][112]=0;ram[73][113]=1;ram[73][114]=1;ram[73][115]=0;ram[73][116]=1;ram[73][117]=1;ram[73][118]=0;ram[73][119]=1;ram[73][120]=0;ram[73][121]=0;ram[73][122]=1;ram[73][123]=0;ram[73][124]=1;ram[73][125]=0;ram[73][126]=0;ram[73][127]=1;ram[73][128]=0;ram[73][129]=0;ram[73][130]=1;ram[73][131]=1;ram[73][132]=0;ram[73][133]=1;ram[73][134]=1;ram[73][135]=1;ram[73][136]=1;
        ram[74][0]=1;ram[74][1]=0;ram[74][2]=1;ram[74][3]=0;ram[74][4]=1;ram[74][5]=1;ram[74][6]=0;ram[74][7]=0;ram[74][8]=1;ram[74][9]=1;ram[74][10]=1;ram[74][11]=1;ram[74][12]=1;ram[74][13]=1;ram[74][14]=0;ram[74][15]=1;ram[74][16]=1;ram[74][17]=0;ram[74][18]=0;ram[74][19]=1;ram[74][20]=0;ram[74][21]=1;ram[74][22]=1;ram[74][23]=1;ram[74][24]=0;ram[74][25]=1;ram[74][26]=1;ram[74][27]=1;ram[74][28]=1;ram[74][29]=0;ram[74][30]=1;ram[74][31]=1;ram[74][32]=0;ram[74][33]=0;ram[74][34]=1;ram[74][35]=0;ram[74][36]=1;ram[74][37]=0;ram[74][38]=1;ram[74][39]=1;ram[74][40]=1;ram[74][41]=0;ram[74][42]=0;ram[74][43]=1;ram[74][44]=0;ram[74][45]=0;ram[74][46]=0;ram[74][47]=0;ram[74][48]=1;ram[74][49]=1;ram[74][50]=0;ram[74][51]=0;ram[74][52]=1;ram[74][53]=0;ram[74][54]=0;ram[74][55]=0;ram[74][56]=1;ram[74][57]=1;ram[74][58]=1;ram[74][59]=1;ram[74][60]=1;ram[74][61]=1;ram[74][62]=1;ram[74][63]=1;ram[74][64]=1;ram[74][65]=1;ram[74][66]=0;ram[74][67]=1;ram[74][68]=1;ram[74][69]=1;ram[74][70]=0;ram[74][71]=0;ram[74][72]=1;ram[74][73]=0;ram[74][74]=0;ram[74][75]=1;ram[74][76]=0;ram[74][77]=1;ram[74][78]=1;ram[74][79]=1;ram[74][80]=1;ram[74][81]=1;ram[74][82]=1;ram[74][83]=1;ram[74][84]=1;ram[74][85]=1;ram[74][86]=1;ram[74][87]=0;ram[74][88]=1;ram[74][89]=0;ram[74][90]=1;ram[74][91]=1;ram[74][92]=1;ram[74][93]=1;ram[74][94]=1;ram[74][95]=0;ram[74][96]=1;ram[74][97]=1;ram[74][98]=0;ram[74][99]=1;ram[74][100]=0;ram[74][101]=0;ram[74][102]=0;ram[74][103]=1;ram[74][104]=0;ram[74][105]=1;ram[74][106]=1;ram[74][107]=1;ram[74][108]=0;ram[74][109]=0;ram[74][110]=1;ram[74][111]=1;ram[74][112]=0;ram[74][113]=1;ram[74][114]=0;ram[74][115]=0;ram[74][116]=1;ram[74][117]=0;ram[74][118]=1;ram[74][119]=1;ram[74][120]=1;ram[74][121]=1;ram[74][122]=0;ram[74][123]=1;ram[74][124]=0;ram[74][125]=1;ram[74][126]=1;ram[74][127]=1;ram[74][128]=1;ram[74][129]=1;ram[74][130]=1;ram[74][131]=1;ram[74][132]=0;ram[74][133]=1;ram[74][134]=1;ram[74][135]=0;ram[74][136]=1;
        ram[75][0]=1;ram[75][1]=1;ram[75][2]=1;ram[75][3]=1;ram[75][4]=0;ram[75][5]=1;ram[75][6]=0;ram[75][7]=0;ram[75][8]=1;ram[75][9]=1;ram[75][10]=1;ram[75][11]=1;ram[75][12]=1;ram[75][13]=1;ram[75][14]=1;ram[75][15]=0;ram[75][16]=1;ram[75][17]=1;ram[75][18]=1;ram[75][19]=0;ram[75][20]=1;ram[75][21]=0;ram[75][22]=1;ram[75][23]=0;ram[75][24]=1;ram[75][25]=1;ram[75][26]=1;ram[75][27]=0;ram[75][28]=0;ram[75][29]=1;ram[75][30]=0;ram[75][31]=1;ram[75][32]=1;ram[75][33]=0;ram[75][34]=1;ram[75][35]=1;ram[75][36]=1;ram[75][37]=1;ram[75][38]=0;ram[75][39]=1;ram[75][40]=0;ram[75][41]=1;ram[75][42]=1;ram[75][43]=1;ram[75][44]=0;ram[75][45]=1;ram[75][46]=1;ram[75][47]=0;ram[75][48]=1;ram[75][49]=1;ram[75][50]=1;ram[75][51]=0;ram[75][52]=1;ram[75][53]=1;ram[75][54]=1;ram[75][55]=1;ram[75][56]=0;ram[75][57]=1;ram[75][58]=0;ram[75][59]=1;ram[75][60]=1;ram[75][61]=0;ram[75][62]=1;ram[75][63]=0;ram[75][64]=0;ram[75][65]=1;ram[75][66]=1;ram[75][67]=1;ram[75][68]=1;ram[75][69]=0;ram[75][70]=1;ram[75][71]=1;ram[75][72]=1;ram[75][73]=1;ram[75][74]=1;ram[75][75]=1;ram[75][76]=1;ram[75][77]=0;ram[75][78]=0;ram[75][79]=1;ram[75][80]=1;ram[75][81]=0;ram[75][82]=1;ram[75][83]=1;ram[75][84]=1;ram[75][85]=1;ram[75][86]=1;ram[75][87]=0;ram[75][88]=1;ram[75][89]=1;ram[75][90]=1;ram[75][91]=0;ram[75][92]=0;ram[75][93]=0;ram[75][94]=1;ram[75][95]=0;ram[75][96]=1;ram[75][97]=0;ram[75][98]=0;ram[75][99]=0;ram[75][100]=0;ram[75][101]=1;ram[75][102]=1;ram[75][103]=1;ram[75][104]=0;ram[75][105]=0;ram[75][106]=0;ram[75][107]=0;ram[75][108]=0;ram[75][109]=1;ram[75][110]=1;ram[75][111]=1;ram[75][112]=1;ram[75][113]=1;ram[75][114]=1;ram[75][115]=1;ram[75][116]=1;ram[75][117]=0;ram[75][118]=1;ram[75][119]=1;ram[75][120]=1;ram[75][121]=1;ram[75][122]=0;ram[75][123]=0;ram[75][124]=0;ram[75][125]=1;ram[75][126]=1;ram[75][127]=0;ram[75][128]=0;ram[75][129]=1;ram[75][130]=1;ram[75][131]=0;ram[75][132]=1;ram[75][133]=0;ram[75][134]=1;ram[75][135]=1;ram[75][136]=1;
        ram[76][0]=0;ram[76][1]=1;ram[76][2]=0;ram[76][3]=1;ram[76][4]=0;ram[76][5]=0;ram[76][6]=1;ram[76][7]=1;ram[76][8]=0;ram[76][9]=1;ram[76][10]=0;ram[76][11]=1;ram[76][12]=1;ram[76][13]=1;ram[76][14]=0;ram[76][15]=0;ram[76][16]=1;ram[76][17]=1;ram[76][18]=1;ram[76][19]=0;ram[76][20]=0;ram[76][21]=1;ram[76][22]=1;ram[76][23]=1;ram[76][24]=1;ram[76][25]=1;ram[76][26]=1;ram[76][27]=1;ram[76][28]=0;ram[76][29]=0;ram[76][30]=1;ram[76][31]=1;ram[76][32]=0;ram[76][33]=0;ram[76][34]=0;ram[76][35]=0;ram[76][36]=1;ram[76][37]=1;ram[76][38]=1;ram[76][39]=0;ram[76][40]=1;ram[76][41]=1;ram[76][42]=0;ram[76][43]=1;ram[76][44]=1;ram[76][45]=1;ram[76][46]=0;ram[76][47]=1;ram[76][48]=1;ram[76][49]=1;ram[76][50]=0;ram[76][51]=1;ram[76][52]=0;ram[76][53]=1;ram[76][54]=1;ram[76][55]=0;ram[76][56]=1;ram[76][57]=1;ram[76][58]=1;ram[76][59]=1;ram[76][60]=1;ram[76][61]=1;ram[76][62]=1;ram[76][63]=1;ram[76][64]=1;ram[76][65]=1;ram[76][66]=1;ram[76][67]=1;ram[76][68]=1;ram[76][69]=1;ram[76][70]=1;ram[76][71]=1;ram[76][72]=1;ram[76][73]=1;ram[76][74]=1;ram[76][75]=1;ram[76][76]=1;ram[76][77]=1;ram[76][78]=1;ram[76][79]=1;ram[76][80]=1;ram[76][81]=0;ram[76][82]=1;ram[76][83]=0;ram[76][84]=1;ram[76][85]=1;ram[76][86]=1;ram[76][87]=1;ram[76][88]=1;ram[76][89]=1;ram[76][90]=1;ram[76][91]=1;ram[76][92]=1;ram[76][93]=1;ram[76][94]=1;ram[76][95]=1;ram[76][96]=0;ram[76][97]=1;ram[76][98]=1;ram[76][99]=1;ram[76][100]=0;ram[76][101]=1;ram[76][102]=0;ram[76][103]=1;ram[76][104]=1;ram[76][105]=0;ram[76][106]=1;ram[76][107]=1;ram[76][108]=1;ram[76][109]=1;ram[76][110]=1;ram[76][111]=1;ram[76][112]=1;ram[76][113]=1;ram[76][114]=1;ram[76][115]=0;ram[76][116]=1;ram[76][117]=1;ram[76][118]=0;ram[76][119]=1;ram[76][120]=1;ram[76][121]=1;ram[76][122]=1;ram[76][123]=0;ram[76][124]=1;ram[76][125]=1;ram[76][126]=0;ram[76][127]=1;ram[76][128]=0;ram[76][129]=1;ram[76][130]=0;ram[76][131]=1;ram[76][132]=1;ram[76][133]=1;ram[76][134]=1;ram[76][135]=1;ram[76][136]=1;
        ram[77][0]=1;ram[77][1]=1;ram[77][2]=1;ram[77][3]=0;ram[77][4]=0;ram[77][5]=1;ram[77][6]=1;ram[77][7]=0;ram[77][8]=1;ram[77][9]=1;ram[77][10]=0;ram[77][11]=1;ram[77][12]=0;ram[77][13]=1;ram[77][14]=1;ram[77][15]=1;ram[77][16]=0;ram[77][17]=1;ram[77][18]=1;ram[77][19]=0;ram[77][20]=0;ram[77][21]=1;ram[77][22]=1;ram[77][23]=0;ram[77][24]=1;ram[77][25]=0;ram[77][26]=0;ram[77][27]=1;ram[77][28]=1;ram[77][29]=0;ram[77][30]=0;ram[77][31]=1;ram[77][32]=1;ram[77][33]=0;ram[77][34]=0;ram[77][35]=1;ram[77][36]=0;ram[77][37]=1;ram[77][38]=1;ram[77][39]=1;ram[77][40]=1;ram[77][41]=1;ram[77][42]=1;ram[77][43]=1;ram[77][44]=1;ram[77][45]=1;ram[77][46]=0;ram[77][47]=1;ram[77][48]=1;ram[77][49]=0;ram[77][50]=1;ram[77][51]=1;ram[77][52]=1;ram[77][53]=1;ram[77][54]=1;ram[77][55]=1;ram[77][56]=0;ram[77][57]=1;ram[77][58]=1;ram[77][59]=1;ram[77][60]=1;ram[77][61]=0;ram[77][62]=1;ram[77][63]=0;ram[77][64]=1;ram[77][65]=1;ram[77][66]=0;ram[77][67]=1;ram[77][68]=0;ram[77][69]=1;ram[77][70]=1;ram[77][71]=1;ram[77][72]=1;ram[77][73]=0;ram[77][74]=0;ram[77][75]=1;ram[77][76]=1;ram[77][77]=1;ram[77][78]=1;ram[77][79]=0;ram[77][80]=1;ram[77][81]=1;ram[77][82]=1;ram[77][83]=0;ram[77][84]=1;ram[77][85]=1;ram[77][86]=1;ram[77][87]=1;ram[77][88]=1;ram[77][89]=1;ram[77][90]=1;ram[77][91]=0;ram[77][92]=1;ram[77][93]=1;ram[77][94]=1;ram[77][95]=1;ram[77][96]=1;ram[77][97]=1;ram[77][98]=0;ram[77][99]=1;ram[77][100]=1;ram[77][101]=1;ram[77][102]=0;ram[77][103]=1;ram[77][104]=1;ram[77][105]=0;ram[77][106]=0;ram[77][107]=1;ram[77][108]=1;ram[77][109]=1;ram[77][110]=1;ram[77][111]=0;ram[77][112]=0;ram[77][113]=1;ram[77][114]=1;ram[77][115]=0;ram[77][116]=0;ram[77][117]=1;ram[77][118]=1;ram[77][119]=1;ram[77][120]=0;ram[77][121]=0;ram[77][122]=0;ram[77][123]=1;ram[77][124]=1;ram[77][125]=1;ram[77][126]=1;ram[77][127]=0;ram[77][128]=0;ram[77][129]=1;ram[77][130]=1;ram[77][131]=0;ram[77][132]=0;ram[77][133]=0;ram[77][134]=0;ram[77][135]=0;ram[77][136]=1;
        ram[78][0]=1;ram[78][1]=0;ram[78][2]=1;ram[78][3]=1;ram[78][4]=1;ram[78][5]=1;ram[78][6]=1;ram[78][7]=0;ram[78][8]=0;ram[78][9]=0;ram[78][10]=1;ram[78][11]=1;ram[78][12]=1;ram[78][13]=0;ram[78][14]=0;ram[78][15]=1;ram[78][16]=1;ram[78][17]=0;ram[78][18]=1;ram[78][19]=0;ram[78][20]=1;ram[78][21]=1;ram[78][22]=1;ram[78][23]=0;ram[78][24]=1;ram[78][25]=0;ram[78][26]=1;ram[78][27]=1;ram[78][28]=0;ram[78][29]=0;ram[78][30]=1;ram[78][31]=1;ram[78][32]=0;ram[78][33]=1;ram[78][34]=0;ram[78][35]=1;ram[78][36]=1;ram[78][37]=1;ram[78][38]=1;ram[78][39]=1;ram[78][40]=1;ram[78][41]=0;ram[78][42]=0;ram[78][43]=0;ram[78][44]=0;ram[78][45]=1;ram[78][46]=1;ram[78][47]=0;ram[78][48]=1;ram[78][49]=0;ram[78][50]=1;ram[78][51]=0;ram[78][52]=1;ram[78][53]=1;ram[78][54]=1;ram[78][55]=1;ram[78][56]=0;ram[78][57]=1;ram[78][58]=1;ram[78][59]=0;ram[78][60]=1;ram[78][61]=1;ram[78][62]=1;ram[78][63]=1;ram[78][64]=1;ram[78][65]=1;ram[78][66]=1;ram[78][67]=1;ram[78][68]=0;ram[78][69]=1;ram[78][70]=0;ram[78][71]=0;ram[78][72]=0;ram[78][73]=1;ram[78][74]=1;ram[78][75]=1;ram[78][76]=0;ram[78][77]=0;ram[78][78]=1;ram[78][79]=1;ram[78][80]=0;ram[78][81]=0;ram[78][82]=1;ram[78][83]=0;ram[78][84]=1;ram[78][85]=1;ram[78][86]=1;ram[78][87]=1;ram[78][88]=1;ram[78][89]=1;ram[78][90]=0;ram[78][91]=1;ram[78][92]=0;ram[78][93]=0;ram[78][94]=1;ram[78][95]=0;ram[78][96]=1;ram[78][97]=1;ram[78][98]=0;ram[78][99]=1;ram[78][100]=1;ram[78][101]=1;ram[78][102]=1;ram[78][103]=1;ram[78][104]=1;ram[78][105]=1;ram[78][106]=1;ram[78][107]=1;ram[78][108]=0;ram[78][109]=0;ram[78][110]=0;ram[78][111]=1;ram[78][112]=1;ram[78][113]=0;ram[78][114]=1;ram[78][115]=1;ram[78][116]=1;ram[78][117]=1;ram[78][118]=1;ram[78][119]=1;ram[78][120]=1;ram[78][121]=0;ram[78][122]=1;ram[78][123]=1;ram[78][124]=0;ram[78][125]=0;ram[78][126]=0;ram[78][127]=1;ram[78][128]=0;ram[78][129]=1;ram[78][130]=1;ram[78][131]=0;ram[78][132]=1;ram[78][133]=1;ram[78][134]=1;ram[78][135]=1;ram[78][136]=1;
        ram[79][0]=1;ram[79][1]=1;ram[79][2]=1;ram[79][3]=1;ram[79][4]=0;ram[79][5]=1;ram[79][6]=1;ram[79][7]=1;ram[79][8]=0;ram[79][9]=1;ram[79][10]=0;ram[79][11]=0;ram[79][12]=0;ram[79][13]=1;ram[79][14]=1;ram[79][15]=0;ram[79][16]=1;ram[79][17]=1;ram[79][18]=1;ram[79][19]=0;ram[79][20]=0;ram[79][21]=1;ram[79][22]=0;ram[79][23]=1;ram[79][24]=1;ram[79][25]=1;ram[79][26]=0;ram[79][27]=1;ram[79][28]=1;ram[79][29]=1;ram[79][30]=1;ram[79][31]=0;ram[79][32]=0;ram[79][33]=1;ram[79][34]=0;ram[79][35]=1;ram[79][36]=1;ram[79][37]=0;ram[79][38]=1;ram[79][39]=1;ram[79][40]=0;ram[79][41]=0;ram[79][42]=1;ram[79][43]=0;ram[79][44]=1;ram[79][45]=1;ram[79][46]=1;ram[79][47]=0;ram[79][48]=1;ram[79][49]=1;ram[79][50]=1;ram[79][51]=1;ram[79][52]=1;ram[79][53]=1;ram[79][54]=0;ram[79][55]=0;ram[79][56]=1;ram[79][57]=1;ram[79][58]=1;ram[79][59]=1;ram[79][60]=1;ram[79][61]=0;ram[79][62]=0;ram[79][63]=1;ram[79][64]=1;ram[79][65]=1;ram[79][66]=0;ram[79][67]=1;ram[79][68]=1;ram[79][69]=0;ram[79][70]=0;ram[79][71]=1;ram[79][72]=1;ram[79][73]=0;ram[79][74]=0;ram[79][75]=1;ram[79][76]=1;ram[79][77]=1;ram[79][78]=1;ram[79][79]=1;ram[79][80]=1;ram[79][81]=1;ram[79][82]=1;ram[79][83]=1;ram[79][84]=1;ram[79][85]=0;ram[79][86]=1;ram[79][87]=0;ram[79][88]=1;ram[79][89]=1;ram[79][90]=0;ram[79][91]=1;ram[79][92]=0;ram[79][93]=0;ram[79][94]=1;ram[79][95]=1;ram[79][96]=1;ram[79][97]=1;ram[79][98]=1;ram[79][99]=1;ram[79][100]=0;ram[79][101]=1;ram[79][102]=1;ram[79][103]=1;ram[79][104]=1;ram[79][105]=1;ram[79][106]=0;ram[79][107]=1;ram[79][108]=1;ram[79][109]=0;ram[79][110]=1;ram[79][111]=1;ram[79][112]=0;ram[79][113]=0;ram[79][114]=1;ram[79][115]=1;ram[79][116]=0;ram[79][117]=1;ram[79][118]=0;ram[79][119]=0;ram[79][120]=0;ram[79][121]=1;ram[79][122]=1;ram[79][123]=1;ram[79][124]=0;ram[79][125]=1;ram[79][126]=1;ram[79][127]=1;ram[79][128]=1;ram[79][129]=1;ram[79][130]=1;ram[79][131]=0;ram[79][132]=1;ram[79][133]=1;ram[79][134]=1;ram[79][135]=1;ram[79][136]=0;
        ram[80][0]=0;ram[80][1]=1;ram[80][2]=1;ram[80][3]=1;ram[80][4]=0;ram[80][5]=0;ram[80][6]=1;ram[80][7]=0;ram[80][8]=1;ram[80][9]=1;ram[80][10]=0;ram[80][11]=0;ram[80][12]=0;ram[80][13]=0;ram[80][14]=0;ram[80][15]=1;ram[80][16]=1;ram[80][17]=1;ram[80][18]=1;ram[80][19]=1;ram[80][20]=1;ram[80][21]=1;ram[80][22]=1;ram[80][23]=1;ram[80][24]=1;ram[80][25]=0;ram[80][26]=1;ram[80][27]=1;ram[80][28]=1;ram[80][29]=1;ram[80][30]=1;ram[80][31]=0;ram[80][32]=1;ram[80][33]=1;ram[80][34]=1;ram[80][35]=1;ram[80][36]=1;ram[80][37]=1;ram[80][38]=0;ram[80][39]=0;ram[80][40]=1;ram[80][41]=0;ram[80][42]=1;ram[80][43]=1;ram[80][44]=1;ram[80][45]=0;ram[80][46]=0;ram[80][47]=0;ram[80][48]=0;ram[80][49]=1;ram[80][50]=1;ram[80][51]=1;ram[80][52]=1;ram[80][53]=1;ram[80][54]=0;ram[80][55]=1;ram[80][56]=0;ram[80][57]=1;ram[80][58]=0;ram[80][59]=1;ram[80][60]=1;ram[80][61]=1;ram[80][62]=1;ram[80][63]=0;ram[80][64]=0;ram[80][65]=0;ram[80][66]=1;ram[80][67]=0;ram[80][68]=1;ram[80][69]=1;ram[80][70]=1;ram[80][71]=1;ram[80][72]=0;ram[80][73]=1;ram[80][74]=1;ram[80][75]=1;ram[80][76]=1;ram[80][77]=1;ram[80][78]=1;ram[80][79]=0;ram[80][80]=1;ram[80][81]=0;ram[80][82]=1;ram[80][83]=1;ram[80][84]=1;ram[80][85]=1;ram[80][86]=0;ram[80][87]=1;ram[80][88]=1;ram[80][89]=1;ram[80][90]=1;ram[80][91]=1;ram[80][92]=1;ram[80][93]=0;ram[80][94]=0;ram[80][95]=0;ram[80][96]=0;ram[80][97]=0;ram[80][98]=0;ram[80][99]=0;ram[80][100]=1;ram[80][101]=0;ram[80][102]=0;ram[80][103]=0;ram[80][104]=0;ram[80][105]=0;ram[80][106]=1;ram[80][107]=1;ram[80][108]=1;ram[80][109]=1;ram[80][110]=1;ram[80][111]=0;ram[80][112]=0;ram[80][113]=0;ram[80][114]=0;ram[80][115]=0;ram[80][116]=1;ram[80][117]=1;ram[80][118]=0;ram[80][119]=1;ram[80][120]=1;ram[80][121]=0;ram[80][122]=1;ram[80][123]=0;ram[80][124]=1;ram[80][125]=1;ram[80][126]=1;ram[80][127]=1;ram[80][128]=0;ram[80][129]=1;ram[80][130]=1;ram[80][131]=0;ram[80][132]=0;ram[80][133]=0;ram[80][134]=0;ram[80][135]=1;ram[80][136]=1;
        ram[81][0]=0;ram[81][1]=1;ram[81][2]=1;ram[81][3]=1;ram[81][4]=1;ram[81][5]=0;ram[81][6]=0;ram[81][7]=1;ram[81][8]=0;ram[81][9]=1;ram[81][10]=1;ram[81][11]=1;ram[81][12]=1;ram[81][13]=0;ram[81][14]=0;ram[81][15]=0;ram[81][16]=1;ram[81][17]=0;ram[81][18]=1;ram[81][19]=0;ram[81][20]=1;ram[81][21]=0;ram[81][22]=0;ram[81][23]=1;ram[81][24]=1;ram[81][25]=1;ram[81][26]=0;ram[81][27]=0;ram[81][28]=1;ram[81][29]=1;ram[81][30]=0;ram[81][31]=1;ram[81][32]=1;ram[81][33]=1;ram[81][34]=0;ram[81][35]=1;ram[81][36]=1;ram[81][37]=0;ram[81][38]=1;ram[81][39]=1;ram[81][40]=0;ram[81][41]=1;ram[81][42]=0;ram[81][43]=1;ram[81][44]=0;ram[81][45]=0;ram[81][46]=0;ram[81][47]=1;ram[81][48]=0;ram[81][49]=0;ram[81][50]=1;ram[81][51]=0;ram[81][52]=1;ram[81][53]=0;ram[81][54]=1;ram[81][55]=1;ram[81][56]=1;ram[81][57]=1;ram[81][58]=1;ram[81][59]=0;ram[81][60]=1;ram[81][61]=1;ram[81][62]=1;ram[81][63]=1;ram[81][64]=1;ram[81][65]=0;ram[81][66]=1;ram[81][67]=1;ram[81][68]=1;ram[81][69]=0;ram[81][70]=1;ram[81][71]=0;ram[81][72]=1;ram[81][73]=1;ram[81][74]=1;ram[81][75]=0;ram[81][76]=1;ram[81][77]=1;ram[81][78]=1;ram[81][79]=0;ram[81][80]=1;ram[81][81]=1;ram[81][82]=1;ram[81][83]=0;ram[81][84]=1;ram[81][85]=0;ram[81][86]=1;ram[81][87]=1;ram[81][88]=1;ram[81][89]=1;ram[81][90]=0;ram[81][91]=0;ram[81][92]=1;ram[81][93]=1;ram[81][94]=0;ram[81][95]=0;ram[81][96]=1;ram[81][97]=1;ram[81][98]=1;ram[81][99]=0;ram[81][100]=0;ram[81][101]=1;ram[81][102]=1;ram[81][103]=0;ram[81][104]=1;ram[81][105]=1;ram[81][106]=0;ram[81][107]=0;ram[81][108]=1;ram[81][109]=1;ram[81][110]=0;ram[81][111]=1;ram[81][112]=1;ram[81][113]=1;ram[81][114]=1;ram[81][115]=0;ram[81][116]=1;ram[81][117]=1;ram[81][118]=0;ram[81][119]=1;ram[81][120]=1;ram[81][121]=1;ram[81][122]=1;ram[81][123]=1;ram[81][124]=1;ram[81][125]=1;ram[81][126]=1;ram[81][127]=1;ram[81][128]=0;ram[81][129]=0;ram[81][130]=0;ram[81][131]=1;ram[81][132]=1;ram[81][133]=1;ram[81][134]=0;ram[81][135]=1;ram[81][136]=1;
        ram[82][0]=0;ram[82][1]=1;ram[82][2]=1;ram[82][3]=1;ram[82][4]=0;ram[82][5]=1;ram[82][6]=1;ram[82][7]=0;ram[82][8]=1;ram[82][9]=1;ram[82][10]=1;ram[82][11]=1;ram[82][12]=1;ram[82][13]=1;ram[82][14]=0;ram[82][15]=0;ram[82][16]=0;ram[82][17]=0;ram[82][18]=0;ram[82][19]=1;ram[82][20]=0;ram[82][21]=0;ram[82][22]=0;ram[82][23]=0;ram[82][24]=1;ram[82][25]=1;ram[82][26]=1;ram[82][27]=0;ram[82][28]=1;ram[82][29]=1;ram[82][30]=0;ram[82][31]=0;ram[82][32]=0;ram[82][33]=0;ram[82][34]=1;ram[82][35]=1;ram[82][36]=0;ram[82][37]=1;ram[82][38]=1;ram[82][39]=1;ram[82][40]=1;ram[82][41]=1;ram[82][42]=1;ram[82][43]=0;ram[82][44]=0;ram[82][45]=1;ram[82][46]=1;ram[82][47]=0;ram[82][48]=1;ram[82][49]=1;ram[82][50]=1;ram[82][51]=1;ram[82][52]=1;ram[82][53]=1;ram[82][54]=1;ram[82][55]=1;ram[82][56]=1;ram[82][57]=1;ram[82][58]=1;ram[82][59]=1;ram[82][60]=0;ram[82][61]=1;ram[82][62]=1;ram[82][63]=1;ram[82][64]=0;ram[82][65]=1;ram[82][66]=0;ram[82][67]=0;ram[82][68]=1;ram[82][69]=1;ram[82][70]=0;ram[82][71]=1;ram[82][72]=1;ram[82][73]=1;ram[82][74]=1;ram[82][75]=1;ram[82][76]=0;ram[82][77]=1;ram[82][78]=1;ram[82][79]=1;ram[82][80]=1;ram[82][81]=1;ram[82][82]=0;ram[82][83]=0;ram[82][84]=0;ram[82][85]=0;ram[82][86]=1;ram[82][87]=1;ram[82][88]=0;ram[82][89]=1;ram[82][90]=1;ram[82][91]=0;ram[82][92]=1;ram[82][93]=1;ram[82][94]=1;ram[82][95]=0;ram[82][96]=1;ram[82][97]=1;ram[82][98]=1;ram[82][99]=0;ram[82][100]=1;ram[82][101]=0;ram[82][102]=0;ram[82][103]=0;ram[82][104]=1;ram[82][105]=1;ram[82][106]=1;ram[82][107]=1;ram[82][108]=1;ram[82][109]=1;ram[82][110]=0;ram[82][111]=1;ram[82][112]=0;ram[82][113]=0;ram[82][114]=1;ram[82][115]=1;ram[82][116]=1;ram[82][117]=1;ram[82][118]=1;ram[82][119]=1;ram[82][120]=0;ram[82][121]=0;ram[82][122]=0;ram[82][123]=1;ram[82][124]=0;ram[82][125]=1;ram[82][126]=0;ram[82][127]=0;ram[82][128]=1;ram[82][129]=1;ram[82][130]=1;ram[82][131]=0;ram[82][132]=1;ram[82][133]=1;ram[82][134]=1;ram[82][135]=0;ram[82][136]=1;
        ram[83][0]=0;ram[83][1]=1;ram[83][2]=1;ram[83][3]=1;ram[83][4]=0;ram[83][5]=0;ram[83][6]=1;ram[83][7]=0;ram[83][8]=1;ram[83][9]=1;ram[83][10]=1;ram[83][11]=0;ram[83][12]=0;ram[83][13]=0;ram[83][14]=1;ram[83][15]=0;ram[83][16]=1;ram[83][17]=1;ram[83][18]=0;ram[83][19]=0;ram[83][20]=0;ram[83][21]=1;ram[83][22]=0;ram[83][23]=1;ram[83][24]=0;ram[83][25]=0;ram[83][26]=1;ram[83][27]=0;ram[83][28]=1;ram[83][29]=0;ram[83][30]=0;ram[83][31]=1;ram[83][32]=0;ram[83][33]=0;ram[83][34]=1;ram[83][35]=0;ram[83][36]=0;ram[83][37]=0;ram[83][38]=0;ram[83][39]=1;ram[83][40]=1;ram[83][41]=1;ram[83][42]=0;ram[83][43]=0;ram[83][44]=0;ram[83][45]=1;ram[83][46]=1;ram[83][47]=1;ram[83][48]=1;ram[83][49]=1;ram[83][50]=1;ram[83][51]=0;ram[83][52]=1;ram[83][53]=0;ram[83][54]=1;ram[83][55]=1;ram[83][56]=0;ram[83][57]=1;ram[83][58]=1;ram[83][59]=1;ram[83][60]=1;ram[83][61]=1;ram[83][62]=1;ram[83][63]=0;ram[83][64]=0;ram[83][65]=1;ram[83][66]=1;ram[83][67]=1;ram[83][68]=1;ram[83][69]=0;ram[83][70]=0;ram[83][71]=1;ram[83][72]=1;ram[83][73]=1;ram[83][74]=1;ram[83][75]=1;ram[83][76]=1;ram[83][77]=1;ram[83][78]=1;ram[83][79]=1;ram[83][80]=0;ram[83][81]=1;ram[83][82]=0;ram[83][83]=0;ram[83][84]=1;ram[83][85]=1;ram[83][86]=1;ram[83][87]=1;ram[83][88]=0;ram[83][89]=0;ram[83][90]=1;ram[83][91]=1;ram[83][92]=1;ram[83][93]=1;ram[83][94]=1;ram[83][95]=1;ram[83][96]=0;ram[83][97]=0;ram[83][98]=1;ram[83][99]=1;ram[83][100]=1;ram[83][101]=0;ram[83][102]=1;ram[83][103]=1;ram[83][104]=0;ram[83][105]=1;ram[83][106]=0;ram[83][107]=1;ram[83][108]=1;ram[83][109]=0;ram[83][110]=1;ram[83][111]=1;ram[83][112]=1;ram[83][113]=0;ram[83][114]=1;ram[83][115]=0;ram[83][116]=0;ram[83][117]=0;ram[83][118]=0;ram[83][119]=0;ram[83][120]=0;ram[83][121]=0;ram[83][122]=1;ram[83][123]=1;ram[83][124]=1;ram[83][125]=1;ram[83][126]=0;ram[83][127]=1;ram[83][128]=0;ram[83][129]=0;ram[83][130]=0;ram[83][131]=1;ram[83][132]=1;ram[83][133]=0;ram[83][134]=0;ram[83][135]=1;ram[83][136]=1;
        ram[84][0]=1;ram[84][1]=1;ram[84][2]=1;ram[84][3]=1;ram[84][4]=0;ram[84][5]=0;ram[84][6]=1;ram[84][7]=1;ram[84][8]=0;ram[84][9]=1;ram[84][10]=0;ram[84][11]=0;ram[84][12]=1;ram[84][13]=0;ram[84][14]=1;ram[84][15]=0;ram[84][16]=1;ram[84][17]=1;ram[84][18]=0;ram[84][19]=1;ram[84][20]=1;ram[84][21]=0;ram[84][22]=0;ram[84][23]=0;ram[84][24]=1;ram[84][25]=0;ram[84][26]=1;ram[84][27]=1;ram[84][28]=0;ram[84][29]=1;ram[84][30]=0;ram[84][31]=0;ram[84][32]=0;ram[84][33]=0;ram[84][34]=1;ram[84][35]=1;ram[84][36]=1;ram[84][37]=1;ram[84][38]=0;ram[84][39]=1;ram[84][40]=0;ram[84][41]=1;ram[84][42]=0;ram[84][43]=1;ram[84][44]=0;ram[84][45]=1;ram[84][46]=0;ram[84][47]=0;ram[84][48]=1;ram[84][49]=0;ram[84][50]=1;ram[84][51]=1;ram[84][52]=1;ram[84][53]=1;ram[84][54]=0;ram[84][55]=0;ram[84][56]=1;ram[84][57]=0;ram[84][58]=1;ram[84][59]=1;ram[84][60]=1;ram[84][61]=1;ram[84][62]=0;ram[84][63]=1;ram[84][64]=1;ram[84][65]=1;ram[84][66]=1;ram[84][67]=1;ram[84][68]=1;ram[84][69]=1;ram[84][70]=1;ram[84][71]=0;ram[84][72]=0;ram[84][73]=1;ram[84][74]=1;ram[84][75]=0;ram[84][76]=0;ram[84][77]=1;ram[84][78]=1;ram[84][79]=1;ram[84][80]=1;ram[84][81]=1;ram[84][82]=1;ram[84][83]=0;ram[84][84]=0;ram[84][85]=1;ram[84][86]=1;ram[84][87]=1;ram[84][88]=0;ram[84][89]=1;ram[84][90]=1;ram[84][91]=1;ram[84][92]=1;ram[84][93]=1;ram[84][94]=0;ram[84][95]=0;ram[84][96]=1;ram[84][97]=1;ram[84][98]=1;ram[84][99]=0;ram[84][100]=1;ram[84][101]=0;ram[84][102]=0;ram[84][103]=1;ram[84][104]=1;ram[84][105]=1;ram[84][106]=1;ram[84][107]=1;ram[84][108]=1;ram[84][109]=0;ram[84][110]=1;ram[84][111]=1;ram[84][112]=0;ram[84][113]=0;ram[84][114]=1;ram[84][115]=1;ram[84][116]=1;ram[84][117]=1;ram[84][118]=0;ram[84][119]=0;ram[84][120]=0;ram[84][121]=1;ram[84][122]=0;ram[84][123]=1;ram[84][124]=1;ram[84][125]=0;ram[84][126]=1;ram[84][127]=0;ram[84][128]=0;ram[84][129]=1;ram[84][130]=0;ram[84][131]=0;ram[84][132]=0;ram[84][133]=0;ram[84][134]=1;ram[84][135]=1;ram[84][136]=0;
        ram[85][0]=1;ram[85][1]=0;ram[85][2]=1;ram[85][3]=1;ram[85][4]=0;ram[85][5]=1;ram[85][6]=0;ram[85][7]=0;ram[85][8]=1;ram[85][9]=1;ram[85][10]=0;ram[85][11]=1;ram[85][12]=0;ram[85][13]=0;ram[85][14]=0;ram[85][15]=0;ram[85][16]=0;ram[85][17]=1;ram[85][18]=1;ram[85][19]=0;ram[85][20]=1;ram[85][21]=1;ram[85][22]=1;ram[85][23]=0;ram[85][24]=1;ram[85][25]=0;ram[85][26]=1;ram[85][27]=0;ram[85][28]=1;ram[85][29]=0;ram[85][30]=1;ram[85][31]=1;ram[85][32]=1;ram[85][33]=1;ram[85][34]=0;ram[85][35]=1;ram[85][36]=1;ram[85][37]=0;ram[85][38]=1;ram[85][39]=1;ram[85][40]=1;ram[85][41]=0;ram[85][42]=0;ram[85][43]=1;ram[85][44]=0;ram[85][45]=0;ram[85][46]=0;ram[85][47]=1;ram[85][48]=1;ram[85][49]=0;ram[85][50]=1;ram[85][51]=1;ram[85][52]=0;ram[85][53]=1;ram[85][54]=0;ram[85][55]=1;ram[85][56]=0;ram[85][57]=0;ram[85][58]=1;ram[85][59]=1;ram[85][60]=1;ram[85][61]=1;ram[85][62]=0;ram[85][63]=0;ram[85][64]=0;ram[85][65]=0;ram[85][66]=0;ram[85][67]=1;ram[85][68]=1;ram[85][69]=1;ram[85][70]=1;ram[85][71]=0;ram[85][72]=0;ram[85][73]=1;ram[85][74]=1;ram[85][75]=1;ram[85][76]=0;ram[85][77]=1;ram[85][78]=0;ram[85][79]=1;ram[85][80]=1;ram[85][81]=0;ram[85][82]=1;ram[85][83]=0;ram[85][84]=1;ram[85][85]=1;ram[85][86]=1;ram[85][87]=0;ram[85][88]=1;ram[85][89]=0;ram[85][90]=1;ram[85][91]=1;ram[85][92]=1;ram[85][93]=0;ram[85][94]=1;ram[85][95]=1;ram[85][96]=1;ram[85][97]=1;ram[85][98]=0;ram[85][99]=1;ram[85][100]=1;ram[85][101]=0;ram[85][102]=1;ram[85][103]=1;ram[85][104]=1;ram[85][105]=1;ram[85][106]=1;ram[85][107]=1;ram[85][108]=0;ram[85][109]=1;ram[85][110]=0;ram[85][111]=1;ram[85][112]=1;ram[85][113]=0;ram[85][114]=1;ram[85][115]=0;ram[85][116]=1;ram[85][117]=1;ram[85][118]=0;ram[85][119]=1;ram[85][120]=1;ram[85][121]=0;ram[85][122]=1;ram[85][123]=1;ram[85][124]=1;ram[85][125]=1;ram[85][126]=0;ram[85][127]=1;ram[85][128]=0;ram[85][129]=0;ram[85][130]=1;ram[85][131]=0;ram[85][132]=0;ram[85][133]=1;ram[85][134]=0;ram[85][135]=1;ram[85][136]=1;
        ram[86][0]=0;ram[86][1]=1;ram[86][2]=0;ram[86][3]=1;ram[86][4]=0;ram[86][5]=0;ram[86][6]=1;ram[86][7]=1;ram[86][8]=1;ram[86][9]=1;ram[86][10]=0;ram[86][11]=1;ram[86][12]=1;ram[86][13]=0;ram[86][14]=0;ram[86][15]=1;ram[86][16]=1;ram[86][17]=1;ram[86][18]=0;ram[86][19]=0;ram[86][20]=0;ram[86][21]=1;ram[86][22]=1;ram[86][23]=1;ram[86][24]=1;ram[86][25]=0;ram[86][26]=0;ram[86][27]=0;ram[86][28]=1;ram[86][29]=1;ram[86][30]=1;ram[86][31]=1;ram[86][32]=0;ram[86][33]=1;ram[86][34]=0;ram[86][35]=0;ram[86][36]=1;ram[86][37]=1;ram[86][38]=1;ram[86][39]=1;ram[86][40]=1;ram[86][41]=1;ram[86][42]=0;ram[86][43]=1;ram[86][44]=0;ram[86][45]=0;ram[86][46]=0;ram[86][47]=1;ram[86][48]=1;ram[86][49]=1;ram[86][50]=0;ram[86][51]=0;ram[86][52]=1;ram[86][53]=0;ram[86][54]=1;ram[86][55]=1;ram[86][56]=0;ram[86][57]=0;ram[86][58]=0;ram[86][59]=1;ram[86][60]=1;ram[86][61]=1;ram[86][62]=0;ram[86][63]=1;ram[86][64]=1;ram[86][65]=1;ram[86][66]=1;ram[86][67]=1;ram[86][68]=0;ram[86][69]=0;ram[86][70]=1;ram[86][71]=1;ram[86][72]=0;ram[86][73]=0;ram[86][74]=0;ram[86][75]=0;ram[86][76]=1;ram[86][77]=1;ram[86][78]=0;ram[86][79]=1;ram[86][80]=1;ram[86][81]=1;ram[86][82]=1;ram[86][83]=1;ram[86][84]=1;ram[86][85]=1;ram[86][86]=1;ram[86][87]=0;ram[86][88]=0;ram[86][89]=1;ram[86][90]=0;ram[86][91]=1;ram[86][92]=0;ram[86][93]=1;ram[86][94]=0;ram[86][95]=1;ram[86][96]=0;ram[86][97]=1;ram[86][98]=1;ram[86][99]=1;ram[86][100]=1;ram[86][101]=0;ram[86][102]=1;ram[86][103]=1;ram[86][104]=1;ram[86][105]=0;ram[86][106]=0;ram[86][107]=1;ram[86][108]=1;ram[86][109]=1;ram[86][110]=1;ram[86][111]=0;ram[86][112]=1;ram[86][113]=1;ram[86][114]=1;ram[86][115]=1;ram[86][116]=1;ram[86][117]=1;ram[86][118]=0;ram[86][119]=0;ram[86][120]=1;ram[86][121]=0;ram[86][122]=1;ram[86][123]=1;ram[86][124]=0;ram[86][125]=1;ram[86][126]=0;ram[86][127]=1;ram[86][128]=1;ram[86][129]=0;ram[86][130]=1;ram[86][131]=1;ram[86][132]=1;ram[86][133]=1;ram[86][134]=0;ram[86][135]=1;ram[86][136]=1;
        ram[87][0]=1;ram[87][1]=0;ram[87][2]=0;ram[87][3]=1;ram[87][4]=1;ram[87][5]=0;ram[87][6]=0;ram[87][7]=0;ram[87][8]=1;ram[87][9]=0;ram[87][10]=1;ram[87][11]=0;ram[87][12]=0;ram[87][13]=0;ram[87][14]=1;ram[87][15]=0;ram[87][16]=0;ram[87][17]=0;ram[87][18]=0;ram[87][19]=1;ram[87][20]=1;ram[87][21]=1;ram[87][22]=1;ram[87][23]=1;ram[87][24]=0;ram[87][25]=1;ram[87][26]=1;ram[87][27]=1;ram[87][28]=0;ram[87][29]=1;ram[87][30]=0;ram[87][31]=0;ram[87][32]=0;ram[87][33]=1;ram[87][34]=0;ram[87][35]=0;ram[87][36]=0;ram[87][37]=1;ram[87][38]=0;ram[87][39]=0;ram[87][40]=1;ram[87][41]=1;ram[87][42]=1;ram[87][43]=0;ram[87][44]=1;ram[87][45]=1;ram[87][46]=1;ram[87][47]=1;ram[87][48]=0;ram[87][49]=0;ram[87][50]=0;ram[87][51]=1;ram[87][52]=1;ram[87][53]=1;ram[87][54]=1;ram[87][55]=1;ram[87][56]=1;ram[87][57]=1;ram[87][58]=0;ram[87][59]=1;ram[87][60]=1;ram[87][61]=1;ram[87][62]=1;ram[87][63]=1;ram[87][64]=1;ram[87][65]=0;ram[87][66]=1;ram[87][67]=1;ram[87][68]=1;ram[87][69]=0;ram[87][70]=1;ram[87][71]=1;ram[87][72]=1;ram[87][73]=1;ram[87][74]=1;ram[87][75]=0;ram[87][76]=1;ram[87][77]=0;ram[87][78]=0;ram[87][79]=0;ram[87][80]=1;ram[87][81]=0;ram[87][82]=0;ram[87][83]=1;ram[87][84]=1;ram[87][85]=1;ram[87][86]=0;ram[87][87]=1;ram[87][88]=0;ram[87][89]=1;ram[87][90]=1;ram[87][91]=0;ram[87][92]=1;ram[87][93]=1;ram[87][94]=1;ram[87][95]=0;ram[87][96]=0;ram[87][97]=1;ram[87][98]=1;ram[87][99]=1;ram[87][100]=1;ram[87][101]=0;ram[87][102]=0;ram[87][103]=0;ram[87][104]=1;ram[87][105]=1;ram[87][106]=0;ram[87][107]=0;ram[87][108]=0;ram[87][109]=1;ram[87][110]=1;ram[87][111]=1;ram[87][112]=0;ram[87][113]=1;ram[87][114]=0;ram[87][115]=0;ram[87][116]=0;ram[87][117]=1;ram[87][118]=1;ram[87][119]=0;ram[87][120]=1;ram[87][121]=1;ram[87][122]=0;ram[87][123]=1;ram[87][124]=0;ram[87][125]=1;ram[87][126]=1;ram[87][127]=0;ram[87][128]=0;ram[87][129]=1;ram[87][130]=0;ram[87][131]=1;ram[87][132]=1;ram[87][133]=1;ram[87][134]=1;ram[87][135]=0;ram[87][136]=0;
        ram[88][0]=1;ram[88][1]=1;ram[88][2]=1;ram[88][3]=1;ram[88][4]=1;ram[88][5]=1;ram[88][6]=1;ram[88][7]=0;ram[88][8]=0;ram[88][9]=0;ram[88][10]=1;ram[88][11]=1;ram[88][12]=1;ram[88][13]=1;ram[88][14]=1;ram[88][15]=0;ram[88][16]=1;ram[88][17]=0;ram[88][18]=0;ram[88][19]=0;ram[88][20]=0;ram[88][21]=1;ram[88][22]=1;ram[88][23]=0;ram[88][24]=1;ram[88][25]=1;ram[88][26]=0;ram[88][27]=0;ram[88][28]=1;ram[88][29]=0;ram[88][30]=1;ram[88][31]=1;ram[88][32]=1;ram[88][33]=1;ram[88][34]=0;ram[88][35]=0;ram[88][36]=1;ram[88][37]=1;ram[88][38]=0;ram[88][39]=0;ram[88][40]=1;ram[88][41]=0;ram[88][42]=0;ram[88][43]=0;ram[88][44]=1;ram[88][45]=1;ram[88][46]=0;ram[88][47]=1;ram[88][48]=1;ram[88][49]=1;ram[88][50]=1;ram[88][51]=1;ram[88][52]=0;ram[88][53]=1;ram[88][54]=1;ram[88][55]=0;ram[88][56]=0;ram[88][57]=1;ram[88][58]=1;ram[88][59]=0;ram[88][60]=0;ram[88][61]=1;ram[88][62]=1;ram[88][63]=1;ram[88][64]=0;ram[88][65]=0;ram[88][66]=1;ram[88][67]=0;ram[88][68]=1;ram[88][69]=1;ram[88][70]=0;ram[88][71]=1;ram[88][72]=0;ram[88][73]=1;ram[88][74]=0;ram[88][75]=0;ram[88][76]=1;ram[88][77]=0;ram[88][78]=0;ram[88][79]=1;ram[88][80]=1;ram[88][81]=0;ram[88][82]=0;ram[88][83]=0;ram[88][84]=1;ram[88][85]=1;ram[88][86]=1;ram[88][87]=0;ram[88][88]=0;ram[88][89]=1;ram[88][90]=0;ram[88][91]=1;ram[88][92]=1;ram[88][93]=1;ram[88][94]=1;ram[88][95]=1;ram[88][96]=0;ram[88][97]=0;ram[88][98]=0;ram[88][99]=1;ram[88][100]=0;ram[88][101]=0;ram[88][102]=1;ram[88][103]=0;ram[88][104]=1;ram[88][105]=1;ram[88][106]=1;ram[88][107]=1;ram[88][108]=1;ram[88][109]=1;ram[88][110]=1;ram[88][111]=1;ram[88][112]=1;ram[88][113]=1;ram[88][114]=0;ram[88][115]=0;ram[88][116]=1;ram[88][117]=0;ram[88][118]=0;ram[88][119]=1;ram[88][120]=0;ram[88][121]=1;ram[88][122]=0;ram[88][123]=1;ram[88][124]=1;ram[88][125]=0;ram[88][126]=1;ram[88][127]=1;ram[88][128]=0;ram[88][129]=1;ram[88][130]=0;ram[88][131]=1;ram[88][132]=0;ram[88][133]=1;ram[88][134]=1;ram[88][135]=0;ram[88][136]=1;
        ram[89][0]=1;ram[89][1]=1;ram[89][2]=1;ram[89][3]=0;ram[89][4]=1;ram[89][5]=1;ram[89][6]=0;ram[89][7]=0;ram[89][8]=1;ram[89][9]=1;ram[89][10]=1;ram[89][11]=0;ram[89][12]=1;ram[89][13]=1;ram[89][14]=1;ram[89][15]=1;ram[89][16]=0;ram[89][17]=1;ram[89][18]=1;ram[89][19]=1;ram[89][20]=1;ram[89][21]=1;ram[89][22]=1;ram[89][23]=0;ram[89][24]=0;ram[89][25]=0;ram[89][26]=1;ram[89][27]=1;ram[89][28]=0;ram[89][29]=0;ram[89][30]=1;ram[89][31]=0;ram[89][32]=1;ram[89][33]=1;ram[89][34]=1;ram[89][35]=1;ram[89][36]=1;ram[89][37]=0;ram[89][38]=0;ram[89][39]=1;ram[89][40]=1;ram[89][41]=1;ram[89][42]=1;ram[89][43]=0;ram[89][44]=0;ram[89][45]=1;ram[89][46]=0;ram[89][47]=1;ram[89][48]=1;ram[89][49]=1;ram[89][50]=1;ram[89][51]=1;ram[89][52]=0;ram[89][53]=1;ram[89][54]=1;ram[89][55]=0;ram[89][56]=0;ram[89][57]=0;ram[89][58]=0;ram[89][59]=0;ram[89][60]=1;ram[89][61]=1;ram[89][62]=1;ram[89][63]=0;ram[89][64]=0;ram[89][65]=1;ram[89][66]=0;ram[89][67]=1;ram[89][68]=1;ram[89][69]=1;ram[89][70]=1;ram[89][71]=0;ram[89][72]=0;ram[89][73]=1;ram[89][74]=0;ram[89][75]=1;ram[89][76]=0;ram[89][77]=0;ram[89][78]=1;ram[89][79]=0;ram[89][80]=1;ram[89][81]=1;ram[89][82]=1;ram[89][83]=1;ram[89][84]=1;ram[89][85]=1;ram[89][86]=0;ram[89][87]=0;ram[89][88]=1;ram[89][89]=1;ram[89][90]=0;ram[89][91]=1;ram[89][92]=1;ram[89][93]=1;ram[89][94]=0;ram[89][95]=1;ram[89][96]=0;ram[89][97]=1;ram[89][98]=0;ram[89][99]=0;ram[89][100]=1;ram[89][101]=1;ram[89][102]=1;ram[89][103]=1;ram[89][104]=1;ram[89][105]=0;ram[89][106]=0;ram[89][107]=0;ram[89][108]=0;ram[89][109]=1;ram[89][110]=0;ram[89][111]=1;ram[89][112]=1;ram[89][113]=1;ram[89][114]=1;ram[89][115]=1;ram[89][116]=1;ram[89][117]=1;ram[89][118]=1;ram[89][119]=0;ram[89][120]=0;ram[89][121]=1;ram[89][122]=0;ram[89][123]=1;ram[89][124]=1;ram[89][125]=1;ram[89][126]=1;ram[89][127]=1;ram[89][128]=0;ram[89][129]=1;ram[89][130]=0;ram[89][131]=1;ram[89][132]=1;ram[89][133]=1;ram[89][134]=1;ram[89][135]=0;ram[89][136]=0;
        ram[90][0]=1;ram[90][1]=1;ram[90][2]=1;ram[90][3]=0;ram[90][4]=1;ram[90][5]=0;ram[90][6]=0;ram[90][7]=0;ram[90][8]=1;ram[90][9]=0;ram[90][10]=1;ram[90][11]=1;ram[90][12]=1;ram[90][13]=1;ram[90][14]=0;ram[90][15]=1;ram[90][16]=0;ram[90][17]=1;ram[90][18]=0;ram[90][19]=1;ram[90][20]=1;ram[90][21]=0;ram[90][22]=1;ram[90][23]=1;ram[90][24]=0;ram[90][25]=1;ram[90][26]=1;ram[90][27]=0;ram[90][28]=0;ram[90][29]=1;ram[90][30]=0;ram[90][31]=1;ram[90][32]=1;ram[90][33]=1;ram[90][34]=1;ram[90][35]=1;ram[90][36]=1;ram[90][37]=1;ram[90][38]=0;ram[90][39]=1;ram[90][40]=1;ram[90][41]=0;ram[90][42]=0;ram[90][43]=1;ram[90][44]=1;ram[90][45]=1;ram[90][46]=0;ram[90][47]=0;ram[90][48]=1;ram[90][49]=1;ram[90][50]=1;ram[90][51]=1;ram[90][52]=0;ram[90][53]=1;ram[90][54]=0;ram[90][55]=0;ram[90][56]=0;ram[90][57]=0;ram[90][58]=1;ram[90][59]=1;ram[90][60]=0;ram[90][61]=1;ram[90][62]=0;ram[90][63]=1;ram[90][64]=1;ram[90][65]=1;ram[90][66]=1;ram[90][67]=1;ram[90][68]=1;ram[90][69]=0;ram[90][70]=1;ram[90][71]=0;ram[90][72]=1;ram[90][73]=1;ram[90][74]=1;ram[90][75]=1;ram[90][76]=1;ram[90][77]=0;ram[90][78]=0;ram[90][79]=1;ram[90][80]=0;ram[90][81]=1;ram[90][82]=1;ram[90][83]=1;ram[90][84]=1;ram[90][85]=1;ram[90][86]=1;ram[90][87]=1;ram[90][88]=0;ram[90][89]=1;ram[90][90]=0;ram[90][91]=1;ram[90][92]=0;ram[90][93]=1;ram[90][94]=1;ram[90][95]=1;ram[90][96]=0;ram[90][97]=0;ram[90][98]=0;ram[90][99]=0;ram[90][100]=1;ram[90][101]=1;ram[90][102]=1;ram[90][103]=0;ram[90][104]=1;ram[90][105]=1;ram[90][106]=1;ram[90][107]=0;ram[90][108]=1;ram[90][109]=1;ram[90][110]=1;ram[90][111]=1;ram[90][112]=0;ram[90][113]=1;ram[90][114]=1;ram[90][115]=0;ram[90][116]=1;ram[90][117]=1;ram[90][118]=1;ram[90][119]=0;ram[90][120]=0;ram[90][121]=1;ram[90][122]=1;ram[90][123]=1;ram[90][124]=1;ram[90][125]=1;ram[90][126]=1;ram[90][127]=1;ram[90][128]=1;ram[90][129]=1;ram[90][130]=1;ram[90][131]=1;ram[90][132]=1;ram[90][133]=1;ram[90][134]=1;ram[90][135]=1;ram[90][136]=1;
        ram[91][0]=1;ram[91][1]=1;ram[91][2]=0;ram[91][3]=0;ram[91][4]=0;ram[91][5]=0;ram[91][6]=0;ram[91][7]=1;ram[91][8]=1;ram[91][9]=0;ram[91][10]=0;ram[91][11]=1;ram[91][12]=0;ram[91][13]=1;ram[91][14]=0;ram[91][15]=0;ram[91][16]=1;ram[91][17]=1;ram[91][18]=1;ram[91][19]=0;ram[91][20]=1;ram[91][21]=0;ram[91][22]=0;ram[91][23]=0;ram[91][24]=1;ram[91][25]=0;ram[91][26]=0;ram[91][27]=0;ram[91][28]=1;ram[91][29]=0;ram[91][30]=0;ram[91][31]=0;ram[91][32]=0;ram[91][33]=1;ram[91][34]=0;ram[91][35]=1;ram[91][36]=1;ram[91][37]=0;ram[91][38]=1;ram[91][39]=0;ram[91][40]=0;ram[91][41]=1;ram[91][42]=0;ram[91][43]=1;ram[91][44]=1;ram[91][45]=0;ram[91][46]=1;ram[91][47]=1;ram[91][48]=1;ram[91][49]=1;ram[91][50]=0;ram[91][51]=1;ram[91][52]=0;ram[91][53]=1;ram[91][54]=0;ram[91][55]=0;ram[91][56]=1;ram[91][57]=0;ram[91][58]=0;ram[91][59]=1;ram[91][60]=0;ram[91][61]=1;ram[91][62]=1;ram[91][63]=1;ram[91][64]=1;ram[91][65]=0;ram[91][66]=1;ram[91][67]=1;ram[91][68]=0;ram[91][69]=0;ram[91][70]=1;ram[91][71]=0;ram[91][72]=1;ram[91][73]=0;ram[91][74]=1;ram[91][75]=0;ram[91][76]=1;ram[91][77]=1;ram[91][78]=0;ram[91][79]=1;ram[91][80]=1;ram[91][81]=1;ram[91][82]=0;ram[91][83]=1;ram[91][84]=0;ram[91][85]=0;ram[91][86]=1;ram[91][87]=1;ram[91][88]=1;ram[91][89]=1;ram[91][90]=1;ram[91][91]=0;ram[91][92]=0;ram[91][93]=1;ram[91][94]=0;ram[91][95]=1;ram[91][96]=0;ram[91][97]=0;ram[91][98]=1;ram[91][99]=0;ram[91][100]=1;ram[91][101]=1;ram[91][102]=0;ram[91][103]=0;ram[91][104]=1;ram[91][105]=0;ram[91][106]=0;ram[91][107]=0;ram[91][108]=0;ram[91][109]=1;ram[91][110]=0;ram[91][111]=1;ram[91][112]=1;ram[91][113]=1;ram[91][114]=0;ram[91][115]=0;ram[91][116]=1;ram[91][117]=0;ram[91][118]=1;ram[91][119]=1;ram[91][120]=0;ram[91][121]=1;ram[91][122]=1;ram[91][123]=1;ram[91][124]=1;ram[91][125]=1;ram[91][126]=1;ram[91][127]=1;ram[91][128]=1;ram[91][129]=0;ram[91][130]=1;ram[91][131]=1;ram[91][132]=1;ram[91][133]=1;ram[91][134]=0;ram[91][135]=1;ram[91][136]=0;
        ram[92][0]=1;ram[92][1]=1;ram[92][2]=1;ram[92][3]=0;ram[92][4]=0;ram[92][5]=0;ram[92][6]=1;ram[92][7]=1;ram[92][8]=1;ram[92][9]=0;ram[92][10]=1;ram[92][11]=0;ram[92][12]=0;ram[92][13]=1;ram[92][14]=0;ram[92][15]=1;ram[92][16]=1;ram[92][17]=0;ram[92][18]=0;ram[92][19]=1;ram[92][20]=0;ram[92][21]=0;ram[92][22]=1;ram[92][23]=0;ram[92][24]=0;ram[92][25]=1;ram[92][26]=1;ram[92][27]=1;ram[92][28]=1;ram[92][29]=0;ram[92][30]=1;ram[92][31]=0;ram[92][32]=1;ram[92][33]=1;ram[92][34]=1;ram[92][35]=0;ram[92][36]=1;ram[92][37]=0;ram[92][38]=1;ram[92][39]=1;ram[92][40]=1;ram[92][41]=1;ram[92][42]=1;ram[92][43]=1;ram[92][44]=1;ram[92][45]=1;ram[92][46]=1;ram[92][47]=0;ram[92][48]=1;ram[92][49]=1;ram[92][50]=1;ram[92][51]=0;ram[92][52]=0;ram[92][53]=1;ram[92][54]=0;ram[92][55]=1;ram[92][56]=1;ram[92][57]=0;ram[92][58]=0;ram[92][59]=1;ram[92][60]=1;ram[92][61]=1;ram[92][62]=1;ram[92][63]=0;ram[92][64]=0;ram[92][65]=1;ram[92][66]=0;ram[92][67]=1;ram[92][68]=0;ram[92][69]=0;ram[92][70]=1;ram[92][71]=1;ram[92][72]=0;ram[92][73]=1;ram[92][74]=1;ram[92][75]=1;ram[92][76]=1;ram[92][77]=1;ram[92][78]=1;ram[92][79]=1;ram[92][80]=0;ram[92][81]=1;ram[92][82]=1;ram[92][83]=1;ram[92][84]=1;ram[92][85]=1;ram[92][86]=1;ram[92][87]=1;ram[92][88]=0;ram[92][89]=1;ram[92][90]=0;ram[92][91]=0;ram[92][92]=1;ram[92][93]=1;ram[92][94]=1;ram[92][95]=0;ram[92][96]=0;ram[92][97]=1;ram[92][98]=1;ram[92][99]=1;ram[92][100]=1;ram[92][101]=1;ram[92][102]=1;ram[92][103]=1;ram[92][104]=0;ram[92][105]=1;ram[92][106]=0;ram[92][107]=0;ram[92][108]=1;ram[92][109]=0;ram[92][110]=1;ram[92][111]=1;ram[92][112]=1;ram[92][113]=1;ram[92][114]=0;ram[92][115]=1;ram[92][116]=1;ram[92][117]=1;ram[92][118]=0;ram[92][119]=0;ram[92][120]=0;ram[92][121]=1;ram[92][122]=1;ram[92][123]=1;ram[92][124]=0;ram[92][125]=1;ram[92][126]=1;ram[92][127]=0;ram[92][128]=1;ram[92][129]=0;ram[92][130]=0;ram[92][131]=1;ram[92][132]=1;ram[92][133]=1;ram[92][134]=0;ram[92][135]=1;ram[92][136]=1;
        ram[93][0]=1;ram[93][1]=1;ram[93][2]=1;ram[93][3]=0;ram[93][4]=1;ram[93][5]=0;ram[93][6]=1;ram[93][7]=0;ram[93][8]=1;ram[93][9]=1;ram[93][10]=1;ram[93][11]=0;ram[93][12]=1;ram[93][13]=0;ram[93][14]=1;ram[93][15]=0;ram[93][16]=0;ram[93][17]=0;ram[93][18]=1;ram[93][19]=1;ram[93][20]=1;ram[93][21]=0;ram[93][22]=0;ram[93][23]=1;ram[93][24]=0;ram[93][25]=0;ram[93][26]=1;ram[93][27]=0;ram[93][28]=1;ram[93][29]=0;ram[93][30]=1;ram[93][31]=1;ram[93][32]=0;ram[93][33]=1;ram[93][34]=1;ram[93][35]=1;ram[93][36]=1;ram[93][37]=1;ram[93][38]=1;ram[93][39]=1;ram[93][40]=1;ram[93][41]=0;ram[93][42]=0;ram[93][43]=1;ram[93][44]=1;ram[93][45]=1;ram[93][46]=1;ram[93][47]=1;ram[93][48]=0;ram[93][49]=1;ram[93][50]=0;ram[93][51]=1;ram[93][52]=0;ram[93][53]=0;ram[93][54]=1;ram[93][55]=1;ram[93][56]=0;ram[93][57]=1;ram[93][58]=0;ram[93][59]=1;ram[93][60]=1;ram[93][61]=0;ram[93][62]=1;ram[93][63]=1;ram[93][64]=1;ram[93][65]=0;ram[93][66]=1;ram[93][67]=0;ram[93][68]=1;ram[93][69]=1;ram[93][70]=0;ram[93][71]=0;ram[93][72]=1;ram[93][73]=0;ram[93][74]=1;ram[93][75]=1;ram[93][76]=1;ram[93][77]=1;ram[93][78]=1;ram[93][79]=1;ram[93][80]=0;ram[93][81]=1;ram[93][82]=0;ram[93][83]=1;ram[93][84]=0;ram[93][85]=1;ram[93][86]=1;ram[93][87]=0;ram[93][88]=0;ram[93][89]=0;ram[93][90]=0;ram[93][91]=0;ram[93][92]=1;ram[93][93]=0;ram[93][94]=0;ram[93][95]=0;ram[93][96]=1;ram[93][97]=1;ram[93][98]=1;ram[93][99]=1;ram[93][100]=1;ram[93][101]=1;ram[93][102]=1;ram[93][103]=1;ram[93][104]=1;ram[93][105]=0;ram[93][106]=1;ram[93][107]=1;ram[93][108]=0;ram[93][109]=1;ram[93][110]=0;ram[93][111]=1;ram[93][112]=0;ram[93][113]=1;ram[93][114]=1;ram[93][115]=1;ram[93][116]=1;ram[93][117]=0;ram[93][118]=1;ram[93][119]=1;ram[93][120]=0;ram[93][121]=1;ram[93][122]=1;ram[93][123]=0;ram[93][124]=1;ram[93][125]=0;ram[93][126]=1;ram[93][127]=1;ram[93][128]=1;ram[93][129]=1;ram[93][130]=1;ram[93][131]=0;ram[93][132]=0;ram[93][133]=0;ram[93][134]=1;ram[93][135]=0;ram[93][136]=1;
        ram[94][0]=1;ram[94][1]=1;ram[94][2]=1;ram[94][3]=0;ram[94][4]=1;ram[94][5]=0;ram[94][6]=1;ram[94][7]=0;ram[94][8]=1;ram[94][9]=1;ram[94][10]=0;ram[94][11]=0;ram[94][12]=1;ram[94][13]=1;ram[94][14]=0;ram[94][15]=1;ram[94][16]=1;ram[94][17]=1;ram[94][18]=1;ram[94][19]=1;ram[94][20]=0;ram[94][21]=1;ram[94][22]=1;ram[94][23]=1;ram[94][24]=1;ram[94][25]=0;ram[94][26]=0;ram[94][27]=1;ram[94][28]=1;ram[94][29]=1;ram[94][30]=1;ram[94][31]=1;ram[94][32]=1;ram[94][33]=1;ram[94][34]=0;ram[94][35]=0;ram[94][36]=0;ram[94][37]=1;ram[94][38]=0;ram[94][39]=0;ram[94][40]=0;ram[94][41]=1;ram[94][42]=0;ram[94][43]=1;ram[94][44]=0;ram[94][45]=1;ram[94][46]=1;ram[94][47]=1;ram[94][48]=0;ram[94][49]=0;ram[94][50]=1;ram[94][51]=1;ram[94][52]=1;ram[94][53]=1;ram[94][54]=1;ram[94][55]=1;ram[94][56]=0;ram[94][57]=1;ram[94][58]=1;ram[94][59]=1;ram[94][60]=1;ram[94][61]=0;ram[94][62]=0;ram[94][63]=1;ram[94][64]=1;ram[94][65]=1;ram[94][66]=0;ram[94][67]=1;ram[94][68]=0;ram[94][69]=0;ram[94][70]=1;ram[94][71]=0;ram[94][72]=1;ram[94][73]=0;ram[94][74]=1;ram[94][75]=1;ram[94][76]=1;ram[94][77]=0;ram[94][78]=1;ram[94][79]=0;ram[94][80]=0;ram[94][81]=1;ram[94][82]=0;ram[94][83]=1;ram[94][84]=1;ram[94][85]=1;ram[94][86]=1;ram[94][87]=1;ram[94][88]=0;ram[94][89]=1;ram[94][90]=1;ram[94][91]=1;ram[94][92]=1;ram[94][93]=0;ram[94][94]=0;ram[94][95]=1;ram[94][96]=1;ram[94][97]=1;ram[94][98]=1;ram[94][99]=0;ram[94][100]=1;ram[94][101]=1;ram[94][102]=1;ram[94][103]=1;ram[94][104]=0;ram[94][105]=0;ram[94][106]=1;ram[94][107]=0;ram[94][108]=1;ram[94][109]=0;ram[94][110]=1;ram[94][111]=0;ram[94][112]=1;ram[94][113]=1;ram[94][114]=1;ram[94][115]=0;ram[94][116]=1;ram[94][117]=1;ram[94][118]=1;ram[94][119]=1;ram[94][120]=0;ram[94][121]=1;ram[94][122]=1;ram[94][123]=1;ram[94][124]=1;ram[94][125]=1;ram[94][126]=1;ram[94][127]=0;ram[94][128]=0;ram[94][129]=1;ram[94][130]=0;ram[94][131]=1;ram[94][132]=1;ram[94][133]=1;ram[94][134]=1;ram[94][135]=0;ram[94][136]=1;
        ram[95][0]=1;ram[95][1]=1;ram[95][2]=1;ram[95][3]=1;ram[95][4]=0;ram[95][5]=1;ram[95][6]=0;ram[95][7]=1;ram[95][8]=1;ram[95][9]=1;ram[95][10]=1;ram[95][11]=1;ram[95][12]=1;ram[95][13]=0;ram[95][14]=1;ram[95][15]=1;ram[95][16]=1;ram[95][17]=1;ram[95][18]=1;ram[95][19]=1;ram[95][20]=0;ram[95][21]=0;ram[95][22]=0;ram[95][23]=0;ram[95][24]=0;ram[95][25]=1;ram[95][26]=0;ram[95][27]=1;ram[95][28]=0;ram[95][29]=1;ram[95][30]=1;ram[95][31]=1;ram[95][32]=0;ram[95][33]=1;ram[95][34]=0;ram[95][35]=1;ram[95][36]=1;ram[95][37]=1;ram[95][38]=1;ram[95][39]=0;ram[95][40]=1;ram[95][41]=1;ram[95][42]=1;ram[95][43]=1;ram[95][44]=1;ram[95][45]=1;ram[95][46]=1;ram[95][47]=0;ram[95][48]=1;ram[95][49]=1;ram[95][50]=0;ram[95][51]=0;ram[95][52]=1;ram[95][53]=1;ram[95][54]=1;ram[95][55]=1;ram[95][56]=1;ram[95][57]=1;ram[95][58]=1;ram[95][59]=1;ram[95][60]=1;ram[95][61]=1;ram[95][62]=1;ram[95][63]=1;ram[95][64]=0;ram[95][65]=0;ram[95][66]=0;ram[95][67]=0;ram[95][68]=1;ram[95][69]=1;ram[95][70]=1;ram[95][71]=1;ram[95][72]=0;ram[95][73]=0;ram[95][74]=0;ram[95][75]=1;ram[95][76]=0;ram[95][77]=1;ram[95][78]=0;ram[95][79]=1;ram[95][80]=0;ram[95][81]=1;ram[95][82]=1;ram[95][83]=0;ram[95][84]=1;ram[95][85]=0;ram[95][86]=1;ram[95][87]=0;ram[95][88]=1;ram[95][89]=0;ram[95][90]=1;ram[95][91]=0;ram[95][92]=0;ram[95][93]=0;ram[95][94]=0;ram[95][95]=0;ram[95][96]=1;ram[95][97]=1;ram[95][98]=0;ram[95][99]=1;ram[95][100]=1;ram[95][101]=1;ram[95][102]=1;ram[95][103]=0;ram[95][104]=1;ram[95][105]=0;ram[95][106]=1;ram[95][107]=1;ram[95][108]=0;ram[95][109]=0;ram[95][110]=0;ram[95][111]=1;ram[95][112]=0;ram[95][113]=0;ram[95][114]=0;ram[95][115]=0;ram[95][116]=1;ram[95][117]=1;ram[95][118]=1;ram[95][119]=1;ram[95][120]=1;ram[95][121]=0;ram[95][122]=0;ram[95][123]=1;ram[95][124]=1;ram[95][125]=0;ram[95][126]=0;ram[95][127]=0;ram[95][128]=1;ram[95][129]=1;ram[95][130]=1;ram[95][131]=1;ram[95][132]=1;ram[95][133]=1;ram[95][134]=0;ram[95][135]=1;ram[95][136]=0;
        ram[96][0]=1;ram[96][1]=0;ram[96][2]=1;ram[96][3]=1;ram[96][4]=1;ram[96][5]=0;ram[96][6]=1;ram[96][7]=1;ram[96][8]=0;ram[96][9]=1;ram[96][10]=1;ram[96][11]=1;ram[96][12]=1;ram[96][13]=0;ram[96][14]=1;ram[96][15]=1;ram[96][16]=0;ram[96][17]=1;ram[96][18]=0;ram[96][19]=0;ram[96][20]=1;ram[96][21]=1;ram[96][22]=0;ram[96][23]=1;ram[96][24]=1;ram[96][25]=1;ram[96][26]=1;ram[96][27]=0;ram[96][28]=0;ram[96][29]=1;ram[96][30]=1;ram[96][31]=1;ram[96][32]=1;ram[96][33]=1;ram[96][34]=1;ram[96][35]=0;ram[96][36]=1;ram[96][37]=0;ram[96][38]=1;ram[96][39]=0;ram[96][40]=0;ram[96][41]=1;ram[96][42]=1;ram[96][43]=1;ram[96][44]=1;ram[96][45]=1;ram[96][46]=1;ram[96][47]=0;ram[96][48]=0;ram[96][49]=1;ram[96][50]=0;ram[96][51]=1;ram[96][52]=0;ram[96][53]=1;ram[96][54]=0;ram[96][55]=1;ram[96][56]=1;ram[96][57]=0;ram[96][58]=1;ram[96][59]=1;ram[96][60]=0;ram[96][61]=0;ram[96][62]=1;ram[96][63]=1;ram[96][64]=1;ram[96][65]=1;ram[96][66]=1;ram[96][67]=0;ram[96][68]=1;ram[96][69]=1;ram[96][70]=1;ram[96][71]=1;ram[96][72]=0;ram[96][73]=0;ram[96][74]=0;ram[96][75]=1;ram[96][76]=1;ram[96][77]=1;ram[96][78]=1;ram[96][79]=1;ram[96][80]=0;ram[96][81]=1;ram[96][82]=1;ram[96][83]=1;ram[96][84]=1;ram[96][85]=0;ram[96][86]=1;ram[96][87]=1;ram[96][88]=1;ram[96][89]=1;ram[96][90]=1;ram[96][91]=1;ram[96][92]=1;ram[96][93]=0;ram[96][94]=0;ram[96][95]=0;ram[96][96]=1;ram[96][97]=0;ram[96][98]=1;ram[96][99]=1;ram[96][100]=0;ram[96][101]=1;ram[96][102]=1;ram[96][103]=1;ram[96][104]=1;ram[96][105]=1;ram[96][106]=0;ram[96][107]=0;ram[96][108]=0;ram[96][109]=1;ram[96][110]=1;ram[96][111]=1;ram[96][112]=1;ram[96][113]=1;ram[96][114]=1;ram[96][115]=1;ram[96][116]=1;ram[96][117]=1;ram[96][118]=1;ram[96][119]=1;ram[96][120]=1;ram[96][121]=0;ram[96][122]=1;ram[96][123]=1;ram[96][124]=1;ram[96][125]=1;ram[96][126]=1;ram[96][127]=0;ram[96][128]=0;ram[96][129]=1;ram[96][130]=0;ram[96][131]=1;ram[96][132]=0;ram[96][133]=0;ram[96][134]=1;ram[96][135]=1;ram[96][136]=1;
        ram[97][0]=0;ram[97][1]=1;ram[97][2]=0;ram[97][3]=0;ram[97][4]=0;ram[97][5]=0;ram[97][6]=0;ram[97][7]=1;ram[97][8]=1;ram[97][9]=0;ram[97][10]=0;ram[97][11]=1;ram[97][12]=1;ram[97][13]=0;ram[97][14]=1;ram[97][15]=0;ram[97][16]=1;ram[97][17]=1;ram[97][18]=1;ram[97][19]=1;ram[97][20]=0;ram[97][21]=1;ram[97][22]=1;ram[97][23]=0;ram[97][24]=1;ram[97][25]=0;ram[97][26]=1;ram[97][27]=1;ram[97][28]=0;ram[97][29]=1;ram[97][30]=1;ram[97][31]=0;ram[97][32]=1;ram[97][33]=0;ram[97][34]=1;ram[97][35]=1;ram[97][36]=1;ram[97][37]=1;ram[97][38]=1;ram[97][39]=0;ram[97][40]=1;ram[97][41]=0;ram[97][42]=1;ram[97][43]=0;ram[97][44]=1;ram[97][45]=1;ram[97][46]=0;ram[97][47]=1;ram[97][48]=0;ram[97][49]=1;ram[97][50]=1;ram[97][51]=1;ram[97][52]=1;ram[97][53]=0;ram[97][54]=1;ram[97][55]=1;ram[97][56]=1;ram[97][57]=1;ram[97][58]=0;ram[97][59]=0;ram[97][60]=0;ram[97][61]=1;ram[97][62]=0;ram[97][63]=1;ram[97][64]=1;ram[97][65]=1;ram[97][66]=1;ram[97][67]=1;ram[97][68]=1;ram[97][69]=1;ram[97][70]=0;ram[97][71]=0;ram[97][72]=1;ram[97][73]=1;ram[97][74]=1;ram[97][75]=0;ram[97][76]=0;ram[97][77]=1;ram[97][78]=1;ram[97][79]=1;ram[97][80]=1;ram[97][81]=1;ram[97][82]=0;ram[97][83]=1;ram[97][84]=1;ram[97][85]=1;ram[97][86]=1;ram[97][87]=0;ram[97][88]=1;ram[97][89]=0;ram[97][90]=1;ram[97][91]=0;ram[97][92]=1;ram[97][93]=0;ram[97][94]=1;ram[97][95]=0;ram[97][96]=0;ram[97][97]=0;ram[97][98]=1;ram[97][99]=0;ram[97][100]=0;ram[97][101]=0;ram[97][102]=1;ram[97][103]=0;ram[97][104]=1;ram[97][105]=1;ram[97][106]=0;ram[97][107]=1;ram[97][108]=1;ram[97][109]=1;ram[97][110]=0;ram[97][111]=0;ram[97][112]=0;ram[97][113]=1;ram[97][114]=1;ram[97][115]=0;ram[97][116]=0;ram[97][117]=1;ram[97][118]=1;ram[97][119]=1;ram[97][120]=0;ram[97][121]=1;ram[97][122]=0;ram[97][123]=1;ram[97][124]=1;ram[97][125]=1;ram[97][126]=1;ram[97][127]=1;ram[97][128]=0;ram[97][129]=1;ram[97][130]=0;ram[97][131]=0;ram[97][132]=1;ram[97][133]=1;ram[97][134]=1;ram[97][135]=0;ram[97][136]=1;
        ram[98][0]=1;ram[98][1]=1;ram[98][2]=1;ram[98][3]=1;ram[98][4]=0;ram[98][5]=1;ram[98][6]=1;ram[98][7]=0;ram[98][8]=0;ram[98][9]=0;ram[98][10]=0;ram[98][11]=0;ram[98][12]=1;ram[98][13]=1;ram[98][14]=0;ram[98][15]=1;ram[98][16]=0;ram[98][17]=1;ram[98][18]=0;ram[98][19]=1;ram[98][20]=1;ram[98][21]=1;ram[98][22]=0;ram[98][23]=1;ram[98][24]=0;ram[98][25]=1;ram[98][26]=0;ram[98][27]=1;ram[98][28]=1;ram[98][29]=1;ram[98][30]=1;ram[98][31]=1;ram[98][32]=0;ram[98][33]=1;ram[98][34]=1;ram[98][35]=1;ram[98][36]=0;ram[98][37]=0;ram[98][38]=0;ram[98][39]=1;ram[98][40]=1;ram[98][41]=1;ram[98][42]=1;ram[98][43]=1;ram[98][44]=1;ram[98][45]=1;ram[98][46]=0;ram[98][47]=1;ram[98][48]=0;ram[98][49]=1;ram[98][50]=1;ram[98][51]=1;ram[98][52]=0;ram[98][53]=1;ram[98][54]=0;ram[98][55]=0;ram[98][56]=0;ram[98][57]=1;ram[98][58]=0;ram[98][59]=1;ram[98][60]=1;ram[98][61]=1;ram[98][62]=1;ram[98][63]=0;ram[98][64]=1;ram[98][65]=1;ram[98][66]=1;ram[98][67]=1;ram[98][68]=1;ram[98][69]=1;ram[98][70]=1;ram[98][71]=1;ram[98][72]=0;ram[98][73]=1;ram[98][74]=1;ram[98][75]=1;ram[98][76]=1;ram[98][77]=1;ram[98][78]=1;ram[98][79]=0;ram[98][80]=0;ram[98][81]=0;ram[98][82]=0;ram[98][83]=1;ram[98][84]=1;ram[98][85]=1;ram[98][86]=1;ram[98][87]=0;ram[98][88]=1;ram[98][89]=1;ram[98][90]=1;ram[98][91]=0;ram[98][92]=0;ram[98][93]=1;ram[98][94]=1;ram[98][95]=0;ram[98][96]=1;ram[98][97]=1;ram[98][98]=1;ram[98][99]=0;ram[98][100]=0;ram[98][101]=1;ram[98][102]=1;ram[98][103]=1;ram[98][104]=1;ram[98][105]=0;ram[98][106]=1;ram[98][107]=1;ram[98][108]=0;ram[98][109]=1;ram[98][110]=1;ram[98][111]=1;ram[98][112]=0;ram[98][113]=0;ram[98][114]=1;ram[98][115]=0;ram[98][116]=1;ram[98][117]=1;ram[98][118]=0;ram[98][119]=1;ram[98][120]=1;ram[98][121]=0;ram[98][122]=1;ram[98][123]=1;ram[98][124]=1;ram[98][125]=1;ram[98][126]=1;ram[98][127]=1;ram[98][128]=1;ram[98][129]=1;ram[98][130]=1;ram[98][131]=1;ram[98][132]=0;ram[98][133]=0;ram[98][134]=1;ram[98][135]=1;ram[98][136]=0;
        ram[99][0]=0;ram[99][1]=1;ram[99][2]=1;ram[99][3]=1;ram[99][4]=1;ram[99][5]=1;ram[99][6]=1;ram[99][7]=1;ram[99][8]=0;ram[99][9]=1;ram[99][10]=1;ram[99][11]=1;ram[99][12]=1;ram[99][13]=0;ram[99][14]=1;ram[99][15]=0;ram[99][16]=1;ram[99][17]=1;ram[99][18]=0;ram[99][19]=0;ram[99][20]=1;ram[99][21]=1;ram[99][22]=1;ram[99][23]=1;ram[99][24]=1;ram[99][25]=1;ram[99][26]=1;ram[99][27]=1;ram[99][28]=1;ram[99][29]=0;ram[99][30]=1;ram[99][31]=1;ram[99][32]=1;ram[99][33]=1;ram[99][34]=1;ram[99][35]=0;ram[99][36]=0;ram[99][37]=0;ram[99][38]=0;ram[99][39]=1;ram[99][40]=0;ram[99][41]=0;ram[99][42]=1;ram[99][43]=0;ram[99][44]=0;ram[99][45]=1;ram[99][46]=1;ram[99][47]=0;ram[99][48]=1;ram[99][49]=1;ram[99][50]=1;ram[99][51]=1;ram[99][52]=1;ram[99][53]=1;ram[99][54]=1;ram[99][55]=0;ram[99][56]=0;ram[99][57]=1;ram[99][58]=0;ram[99][59]=0;ram[99][60]=1;ram[99][61]=1;ram[99][62]=1;ram[99][63]=0;ram[99][64]=0;ram[99][65]=0;ram[99][66]=1;ram[99][67]=1;ram[99][68]=1;ram[99][69]=1;ram[99][70]=1;ram[99][71]=1;ram[99][72]=0;ram[99][73]=1;ram[99][74]=1;ram[99][75]=0;ram[99][76]=1;ram[99][77]=1;ram[99][78]=0;ram[99][79]=0;ram[99][80]=1;ram[99][81]=1;ram[99][82]=1;ram[99][83]=1;ram[99][84]=1;ram[99][85]=0;ram[99][86]=0;ram[99][87]=0;ram[99][88]=1;ram[99][89]=1;ram[99][90]=1;ram[99][91]=1;ram[99][92]=0;ram[99][93]=1;ram[99][94]=1;ram[99][95]=1;ram[99][96]=1;ram[99][97]=0;ram[99][98]=0;ram[99][99]=1;ram[99][100]=0;ram[99][101]=1;ram[99][102]=0;ram[99][103]=1;ram[99][104]=1;ram[99][105]=1;ram[99][106]=1;ram[99][107]=0;ram[99][108]=0;ram[99][109]=1;ram[99][110]=1;ram[99][111]=1;ram[99][112]=1;ram[99][113]=0;ram[99][114]=0;ram[99][115]=1;ram[99][116]=0;ram[99][117]=0;ram[99][118]=0;ram[99][119]=1;ram[99][120]=1;ram[99][121]=0;ram[99][122]=1;ram[99][123]=1;ram[99][124]=1;ram[99][125]=1;ram[99][126]=1;ram[99][127]=1;ram[99][128]=1;ram[99][129]=0;ram[99][130]=1;ram[99][131]=1;ram[99][132]=0;ram[99][133]=0;ram[99][134]=0;ram[99][135]=0;ram[99][136]=0;
        ram[100][0]=1;ram[100][1]=0;ram[100][2]=1;ram[100][3]=0;ram[100][4]=1;ram[100][5]=0;ram[100][6]=1;ram[100][7]=1;ram[100][8]=1;ram[100][9]=1;ram[100][10]=1;ram[100][11]=1;ram[100][12]=1;ram[100][13]=0;ram[100][14]=0;ram[100][15]=0;ram[100][16]=1;ram[100][17]=1;ram[100][18]=0;ram[100][19]=1;ram[100][20]=1;ram[100][21]=1;ram[100][22]=0;ram[100][23]=0;ram[100][24]=0;ram[100][25]=1;ram[100][26]=0;ram[100][27]=1;ram[100][28]=1;ram[100][29]=0;ram[100][30]=1;ram[100][31]=0;ram[100][32]=0;ram[100][33]=1;ram[100][34]=0;ram[100][35]=1;ram[100][36]=0;ram[100][37]=1;ram[100][38]=0;ram[100][39]=1;ram[100][40]=1;ram[100][41]=1;ram[100][42]=0;ram[100][43]=1;ram[100][44]=1;ram[100][45]=0;ram[100][46]=0;ram[100][47]=1;ram[100][48]=1;ram[100][49]=1;ram[100][50]=0;ram[100][51]=1;ram[100][52]=1;ram[100][53]=1;ram[100][54]=1;ram[100][55]=0;ram[100][56]=0;ram[100][57]=1;ram[100][58]=0;ram[100][59]=0;ram[100][60]=0;ram[100][61]=0;ram[100][62]=1;ram[100][63]=0;ram[100][64]=0;ram[100][65]=1;ram[100][66]=1;ram[100][67]=1;ram[100][68]=0;ram[100][69]=1;ram[100][70]=0;ram[100][71]=0;ram[100][72]=1;ram[100][73]=0;ram[100][74]=1;ram[100][75]=0;ram[100][76]=0;ram[100][77]=0;ram[100][78]=0;ram[100][79]=1;ram[100][80]=0;ram[100][81]=1;ram[100][82]=1;ram[100][83]=1;ram[100][84]=0;ram[100][85]=1;ram[100][86]=0;ram[100][87]=1;ram[100][88]=0;ram[100][89]=1;ram[100][90]=1;ram[100][91]=0;ram[100][92]=1;ram[100][93]=1;ram[100][94]=1;ram[100][95]=0;ram[100][96]=1;ram[100][97]=1;ram[100][98]=1;ram[100][99]=1;ram[100][100]=0;ram[100][101]=0;ram[100][102]=1;ram[100][103]=1;ram[100][104]=1;ram[100][105]=1;ram[100][106]=0;ram[100][107]=1;ram[100][108]=1;ram[100][109]=1;ram[100][110]=1;ram[100][111]=0;ram[100][112]=1;ram[100][113]=1;ram[100][114]=1;ram[100][115]=1;ram[100][116]=1;ram[100][117]=1;ram[100][118]=1;ram[100][119]=1;ram[100][120]=1;ram[100][121]=1;ram[100][122]=1;ram[100][123]=1;ram[100][124]=0;ram[100][125]=0;ram[100][126]=1;ram[100][127]=0;ram[100][128]=0;ram[100][129]=0;ram[100][130]=0;ram[100][131]=1;ram[100][132]=1;ram[100][133]=0;ram[100][134]=1;ram[100][135]=1;ram[100][136]=1;
        ram[101][0]=1;ram[101][1]=0;ram[101][2]=1;ram[101][3]=1;ram[101][4]=1;ram[101][5]=0;ram[101][6]=1;ram[101][7]=0;ram[101][8]=1;ram[101][9]=1;ram[101][10]=1;ram[101][11]=1;ram[101][12]=0;ram[101][13]=1;ram[101][14]=1;ram[101][15]=0;ram[101][16]=1;ram[101][17]=1;ram[101][18]=1;ram[101][19]=1;ram[101][20]=1;ram[101][21]=0;ram[101][22]=1;ram[101][23]=1;ram[101][24]=1;ram[101][25]=1;ram[101][26]=1;ram[101][27]=1;ram[101][28]=1;ram[101][29]=1;ram[101][30]=1;ram[101][31]=1;ram[101][32]=1;ram[101][33]=1;ram[101][34]=1;ram[101][35]=1;ram[101][36]=1;ram[101][37]=1;ram[101][38]=0;ram[101][39]=0;ram[101][40]=1;ram[101][41]=0;ram[101][42]=1;ram[101][43]=1;ram[101][44]=1;ram[101][45]=1;ram[101][46]=0;ram[101][47]=1;ram[101][48]=1;ram[101][49]=1;ram[101][50]=1;ram[101][51]=1;ram[101][52]=0;ram[101][53]=0;ram[101][54]=1;ram[101][55]=1;ram[101][56]=1;ram[101][57]=1;ram[101][58]=1;ram[101][59]=1;ram[101][60]=1;ram[101][61]=0;ram[101][62]=1;ram[101][63]=0;ram[101][64]=1;ram[101][65]=1;ram[101][66]=1;ram[101][67]=1;ram[101][68]=0;ram[101][69]=1;ram[101][70]=0;ram[101][71]=1;ram[101][72]=0;ram[101][73]=1;ram[101][74]=1;ram[101][75]=1;ram[101][76]=1;ram[101][77]=1;ram[101][78]=0;ram[101][79]=1;ram[101][80]=1;ram[101][81]=0;ram[101][82]=1;ram[101][83]=0;ram[101][84]=1;ram[101][85]=1;ram[101][86]=1;ram[101][87]=1;ram[101][88]=1;ram[101][89]=0;ram[101][90]=0;ram[101][91]=1;ram[101][92]=1;ram[101][93]=0;ram[101][94]=1;ram[101][95]=0;ram[101][96]=1;ram[101][97]=1;ram[101][98]=1;ram[101][99]=0;ram[101][100]=0;ram[101][101]=1;ram[101][102]=1;ram[101][103]=1;ram[101][104]=1;ram[101][105]=0;ram[101][106]=1;ram[101][107]=1;ram[101][108]=1;ram[101][109]=1;ram[101][110]=0;ram[101][111]=1;ram[101][112]=0;ram[101][113]=0;ram[101][114]=1;ram[101][115]=1;ram[101][116]=0;ram[101][117]=1;ram[101][118]=1;ram[101][119]=0;ram[101][120]=1;ram[101][121]=1;ram[101][122]=1;ram[101][123]=0;ram[101][124]=1;ram[101][125]=0;ram[101][126]=1;ram[101][127]=1;ram[101][128]=0;ram[101][129]=0;ram[101][130]=1;ram[101][131]=1;ram[101][132]=1;ram[101][133]=0;ram[101][134]=0;ram[101][135]=1;ram[101][136]=1;
        ram[102][0]=0;ram[102][1]=1;ram[102][2]=1;ram[102][3]=1;ram[102][4]=1;ram[102][5]=0;ram[102][6]=1;ram[102][7]=1;ram[102][8]=0;ram[102][9]=1;ram[102][10]=1;ram[102][11]=0;ram[102][12]=1;ram[102][13]=1;ram[102][14]=1;ram[102][15]=0;ram[102][16]=1;ram[102][17]=0;ram[102][18]=1;ram[102][19]=0;ram[102][20]=1;ram[102][21]=1;ram[102][22]=1;ram[102][23]=1;ram[102][24]=1;ram[102][25]=0;ram[102][26]=1;ram[102][27]=1;ram[102][28]=1;ram[102][29]=1;ram[102][30]=0;ram[102][31]=0;ram[102][32]=1;ram[102][33]=1;ram[102][34]=1;ram[102][35]=1;ram[102][36]=1;ram[102][37]=1;ram[102][38]=0;ram[102][39]=0;ram[102][40]=1;ram[102][41]=0;ram[102][42]=1;ram[102][43]=1;ram[102][44]=1;ram[102][45]=1;ram[102][46]=0;ram[102][47]=1;ram[102][48]=1;ram[102][49]=0;ram[102][50]=1;ram[102][51]=0;ram[102][52]=1;ram[102][53]=0;ram[102][54]=1;ram[102][55]=1;ram[102][56]=0;ram[102][57]=0;ram[102][58]=1;ram[102][59]=0;ram[102][60]=0;ram[102][61]=1;ram[102][62]=1;ram[102][63]=0;ram[102][64]=0;ram[102][65]=0;ram[102][66]=0;ram[102][67]=1;ram[102][68]=1;ram[102][69]=1;ram[102][70]=1;ram[102][71]=1;ram[102][72]=0;ram[102][73]=1;ram[102][74]=0;ram[102][75]=1;ram[102][76]=0;ram[102][77]=1;ram[102][78]=1;ram[102][79]=0;ram[102][80]=0;ram[102][81]=0;ram[102][82]=1;ram[102][83]=0;ram[102][84]=1;ram[102][85]=1;ram[102][86]=1;ram[102][87]=0;ram[102][88]=0;ram[102][89]=1;ram[102][90]=1;ram[102][91]=0;ram[102][92]=1;ram[102][93]=1;ram[102][94]=1;ram[102][95]=1;ram[102][96]=1;ram[102][97]=1;ram[102][98]=1;ram[102][99]=1;ram[102][100]=0;ram[102][101]=1;ram[102][102]=0;ram[102][103]=1;ram[102][104]=1;ram[102][105]=0;ram[102][106]=0;ram[102][107]=0;ram[102][108]=1;ram[102][109]=0;ram[102][110]=1;ram[102][111]=0;ram[102][112]=0;ram[102][113]=1;ram[102][114]=1;ram[102][115]=0;ram[102][116]=1;ram[102][117]=1;ram[102][118]=1;ram[102][119]=0;ram[102][120]=1;ram[102][121]=1;ram[102][122]=1;ram[102][123]=1;ram[102][124]=1;ram[102][125]=1;ram[102][126]=1;ram[102][127]=1;ram[102][128]=1;ram[102][129]=1;ram[102][130]=1;ram[102][131]=0;ram[102][132]=1;ram[102][133]=1;ram[102][134]=0;ram[102][135]=1;ram[102][136]=1;
        ram[103][0]=1;ram[103][1]=0;ram[103][2]=1;ram[103][3]=1;ram[103][4]=0;ram[103][5]=0;ram[103][6]=0;ram[103][7]=1;ram[103][8]=1;ram[103][9]=1;ram[103][10]=0;ram[103][11]=1;ram[103][12]=1;ram[103][13]=1;ram[103][14]=0;ram[103][15]=1;ram[103][16]=1;ram[103][17]=1;ram[103][18]=1;ram[103][19]=0;ram[103][20]=1;ram[103][21]=1;ram[103][22]=1;ram[103][23]=0;ram[103][24]=0;ram[103][25]=1;ram[103][26]=1;ram[103][27]=0;ram[103][28]=1;ram[103][29]=0;ram[103][30]=1;ram[103][31]=1;ram[103][32]=1;ram[103][33]=1;ram[103][34]=1;ram[103][35]=1;ram[103][36]=1;ram[103][37]=1;ram[103][38]=1;ram[103][39]=1;ram[103][40]=0;ram[103][41]=1;ram[103][42]=1;ram[103][43]=1;ram[103][44]=1;ram[103][45]=1;ram[103][46]=0;ram[103][47]=1;ram[103][48]=1;ram[103][49]=1;ram[103][50]=1;ram[103][51]=1;ram[103][52]=1;ram[103][53]=1;ram[103][54]=0;ram[103][55]=1;ram[103][56]=0;ram[103][57]=0;ram[103][58]=0;ram[103][59]=1;ram[103][60]=1;ram[103][61]=0;ram[103][62]=1;ram[103][63]=0;ram[103][64]=1;ram[103][65]=1;ram[103][66]=1;ram[103][67]=0;ram[103][68]=1;ram[103][69]=0;ram[103][70]=1;ram[103][71]=0;ram[103][72]=1;ram[103][73]=1;ram[103][74]=1;ram[103][75]=1;ram[103][76]=0;ram[103][77]=0;ram[103][78]=1;ram[103][79]=1;ram[103][80]=0;ram[103][81]=1;ram[103][82]=1;ram[103][83]=0;ram[103][84]=1;ram[103][85]=1;ram[103][86]=0;ram[103][87]=1;ram[103][88]=1;ram[103][89]=1;ram[103][90]=1;ram[103][91]=1;ram[103][92]=0;ram[103][93]=0;ram[103][94]=1;ram[103][95]=0;ram[103][96]=1;ram[103][97]=1;ram[103][98]=1;ram[103][99]=0;ram[103][100]=0;ram[103][101]=0;ram[103][102]=0;ram[103][103]=1;ram[103][104]=1;ram[103][105]=1;ram[103][106]=1;ram[103][107]=1;ram[103][108]=1;ram[103][109]=0;ram[103][110]=0;ram[103][111]=0;ram[103][112]=0;ram[103][113]=1;ram[103][114]=1;ram[103][115]=0;ram[103][116]=0;ram[103][117]=1;ram[103][118]=0;ram[103][119]=1;ram[103][120]=1;ram[103][121]=1;ram[103][122]=1;ram[103][123]=1;ram[103][124]=1;ram[103][125]=1;ram[103][126]=1;ram[103][127]=0;ram[103][128]=0;ram[103][129]=1;ram[103][130]=1;ram[103][131]=1;ram[103][132]=1;ram[103][133]=1;ram[103][134]=1;ram[103][135]=1;ram[103][136]=1;
        ram[104][0]=0;ram[104][1]=1;ram[104][2]=0;ram[104][3]=1;ram[104][4]=1;ram[104][5]=0;ram[104][6]=1;ram[104][7]=1;ram[104][8]=0;ram[104][9]=1;ram[104][10]=0;ram[104][11]=0;ram[104][12]=1;ram[104][13]=1;ram[104][14]=1;ram[104][15]=1;ram[104][16]=1;ram[104][17]=1;ram[104][18]=1;ram[104][19]=0;ram[104][20]=1;ram[104][21]=0;ram[104][22]=1;ram[104][23]=1;ram[104][24]=1;ram[104][25]=0;ram[104][26]=0;ram[104][27]=0;ram[104][28]=1;ram[104][29]=0;ram[104][30]=1;ram[104][31]=0;ram[104][32]=1;ram[104][33]=0;ram[104][34]=1;ram[104][35]=1;ram[104][36]=1;ram[104][37]=1;ram[104][38]=1;ram[104][39]=1;ram[104][40]=1;ram[104][41]=1;ram[104][42]=0;ram[104][43]=1;ram[104][44]=1;ram[104][45]=1;ram[104][46]=0;ram[104][47]=1;ram[104][48]=1;ram[104][49]=0;ram[104][50]=1;ram[104][51]=1;ram[104][52]=1;ram[104][53]=1;ram[104][54]=1;ram[104][55]=1;ram[104][56]=1;ram[104][57]=0;ram[104][58]=1;ram[104][59]=0;ram[104][60]=1;ram[104][61]=0;ram[104][62]=1;ram[104][63]=1;ram[104][64]=1;ram[104][65]=0;ram[104][66]=1;ram[104][67]=1;ram[104][68]=1;ram[104][69]=1;ram[104][70]=1;ram[104][71]=1;ram[104][72]=1;ram[104][73]=1;ram[104][74]=0;ram[104][75]=1;ram[104][76]=0;ram[104][77]=1;ram[104][78]=1;ram[104][79]=0;ram[104][80]=0;ram[104][81]=0;ram[104][82]=1;ram[104][83]=1;ram[104][84]=0;ram[104][85]=0;ram[104][86]=1;ram[104][87]=0;ram[104][88]=0;ram[104][89]=1;ram[104][90]=1;ram[104][91]=0;ram[104][92]=1;ram[104][93]=1;ram[104][94]=1;ram[104][95]=1;ram[104][96]=0;ram[104][97]=0;ram[104][98]=1;ram[104][99]=1;ram[104][100]=0;ram[104][101]=1;ram[104][102]=1;ram[104][103]=0;ram[104][104]=1;ram[104][105]=1;ram[104][106]=1;ram[104][107]=0;ram[104][108]=0;ram[104][109]=1;ram[104][110]=0;ram[104][111]=0;ram[104][112]=1;ram[104][113]=1;ram[104][114]=0;ram[104][115]=1;ram[104][116]=1;ram[104][117]=1;ram[104][118]=0;ram[104][119]=1;ram[104][120]=1;ram[104][121]=1;ram[104][122]=1;ram[104][123]=1;ram[104][124]=1;ram[104][125]=1;ram[104][126]=1;ram[104][127]=1;ram[104][128]=1;ram[104][129]=1;ram[104][130]=0;ram[104][131]=1;ram[104][132]=0;ram[104][133]=0;ram[104][134]=1;ram[104][135]=1;ram[104][136]=1;
        ram[105][0]=1;ram[105][1]=1;ram[105][2]=1;ram[105][3]=0;ram[105][4]=0;ram[105][5]=1;ram[105][6]=1;ram[105][7]=1;ram[105][8]=1;ram[105][9]=1;ram[105][10]=1;ram[105][11]=1;ram[105][12]=1;ram[105][13]=1;ram[105][14]=1;ram[105][15]=1;ram[105][16]=1;ram[105][17]=1;ram[105][18]=0;ram[105][19]=0;ram[105][20]=1;ram[105][21]=0;ram[105][22]=1;ram[105][23]=1;ram[105][24]=1;ram[105][25]=0;ram[105][26]=0;ram[105][27]=0;ram[105][28]=1;ram[105][29]=1;ram[105][30]=0;ram[105][31]=1;ram[105][32]=1;ram[105][33]=1;ram[105][34]=1;ram[105][35]=0;ram[105][36]=0;ram[105][37]=1;ram[105][38]=1;ram[105][39]=1;ram[105][40]=1;ram[105][41]=0;ram[105][42]=1;ram[105][43]=1;ram[105][44]=0;ram[105][45]=1;ram[105][46]=1;ram[105][47]=0;ram[105][48]=1;ram[105][49]=1;ram[105][50]=1;ram[105][51]=1;ram[105][52]=1;ram[105][53]=1;ram[105][54]=0;ram[105][55]=0;ram[105][56]=0;ram[105][57]=1;ram[105][58]=0;ram[105][59]=1;ram[105][60]=0;ram[105][61]=1;ram[105][62]=1;ram[105][63]=1;ram[105][64]=1;ram[105][65]=1;ram[105][66]=0;ram[105][67]=1;ram[105][68]=0;ram[105][69]=1;ram[105][70]=1;ram[105][71]=0;ram[105][72]=1;ram[105][73]=0;ram[105][74]=1;ram[105][75]=1;ram[105][76]=1;ram[105][77]=1;ram[105][78]=1;ram[105][79]=0;ram[105][80]=1;ram[105][81]=1;ram[105][82]=1;ram[105][83]=1;ram[105][84]=0;ram[105][85]=0;ram[105][86]=0;ram[105][87]=1;ram[105][88]=0;ram[105][89]=1;ram[105][90]=1;ram[105][91]=1;ram[105][92]=0;ram[105][93]=1;ram[105][94]=0;ram[105][95]=1;ram[105][96]=1;ram[105][97]=0;ram[105][98]=1;ram[105][99]=1;ram[105][100]=1;ram[105][101]=1;ram[105][102]=1;ram[105][103]=0;ram[105][104]=1;ram[105][105]=1;ram[105][106]=1;ram[105][107]=1;ram[105][108]=0;ram[105][109]=1;ram[105][110]=0;ram[105][111]=0;ram[105][112]=1;ram[105][113]=1;ram[105][114]=1;ram[105][115]=0;ram[105][116]=0;ram[105][117]=1;ram[105][118]=0;ram[105][119]=0;ram[105][120]=1;ram[105][121]=1;ram[105][122]=1;ram[105][123]=1;ram[105][124]=0;ram[105][125]=1;ram[105][126]=1;ram[105][127]=0;ram[105][128]=1;ram[105][129]=0;ram[105][130]=0;ram[105][131]=1;ram[105][132]=0;ram[105][133]=1;ram[105][134]=1;ram[105][135]=1;ram[105][136]=0;
        ram[106][0]=1;ram[106][1]=1;ram[106][2]=1;ram[106][3]=1;ram[106][4]=0;ram[106][5]=1;ram[106][6]=1;ram[106][7]=1;ram[106][8]=0;ram[106][9]=1;ram[106][10]=0;ram[106][11]=0;ram[106][12]=0;ram[106][13]=0;ram[106][14]=1;ram[106][15]=1;ram[106][16]=1;ram[106][17]=1;ram[106][18]=1;ram[106][19]=1;ram[106][20]=1;ram[106][21]=0;ram[106][22]=1;ram[106][23]=0;ram[106][24]=0;ram[106][25]=0;ram[106][26]=0;ram[106][27]=1;ram[106][28]=1;ram[106][29]=1;ram[106][30]=0;ram[106][31]=1;ram[106][32]=0;ram[106][33]=0;ram[106][34]=0;ram[106][35]=1;ram[106][36]=1;ram[106][37]=1;ram[106][38]=1;ram[106][39]=1;ram[106][40]=0;ram[106][41]=0;ram[106][42]=0;ram[106][43]=1;ram[106][44]=1;ram[106][45]=1;ram[106][46]=1;ram[106][47]=0;ram[106][48]=1;ram[106][49]=1;ram[106][50]=0;ram[106][51]=1;ram[106][52]=1;ram[106][53]=1;ram[106][54]=1;ram[106][55]=0;ram[106][56]=0;ram[106][57]=0;ram[106][58]=0;ram[106][59]=1;ram[106][60]=0;ram[106][61]=1;ram[106][62]=1;ram[106][63]=1;ram[106][64]=1;ram[106][65]=1;ram[106][66]=0;ram[106][67]=1;ram[106][68]=1;ram[106][69]=0;ram[106][70]=1;ram[106][71]=1;ram[106][72]=1;ram[106][73]=1;ram[106][74]=1;ram[106][75]=1;ram[106][76]=1;ram[106][77]=0;ram[106][78]=0;ram[106][79]=1;ram[106][80]=1;ram[106][81]=0;ram[106][82]=1;ram[106][83]=1;ram[106][84]=0;ram[106][85]=1;ram[106][86]=0;ram[106][87]=1;ram[106][88]=1;ram[106][89]=0;ram[106][90]=1;ram[106][91]=1;ram[106][92]=1;ram[106][93]=0;ram[106][94]=1;ram[106][95]=0;ram[106][96]=1;ram[106][97]=0;ram[106][98]=1;ram[106][99]=1;ram[106][100]=0;ram[106][101]=1;ram[106][102]=0;ram[106][103]=1;ram[106][104]=1;ram[106][105]=1;ram[106][106]=1;ram[106][107]=0;ram[106][108]=1;ram[106][109]=1;ram[106][110]=0;ram[106][111]=0;ram[106][112]=1;ram[106][113]=1;ram[106][114]=1;ram[106][115]=1;ram[106][116]=0;ram[106][117]=1;ram[106][118]=1;ram[106][119]=1;ram[106][120]=1;ram[106][121]=0;ram[106][122]=1;ram[106][123]=1;ram[106][124]=1;ram[106][125]=1;ram[106][126]=1;ram[106][127]=0;ram[106][128]=0;ram[106][129]=1;ram[106][130]=0;ram[106][131]=1;ram[106][132]=0;ram[106][133]=1;ram[106][134]=0;ram[106][135]=0;ram[106][136]=1;
        ram[107][0]=1;ram[107][1]=1;ram[107][2]=0;ram[107][3]=0;ram[107][4]=1;ram[107][5]=1;ram[107][6]=1;ram[107][7]=0;ram[107][8]=0;ram[107][9]=1;ram[107][10]=1;ram[107][11]=0;ram[107][12]=1;ram[107][13]=1;ram[107][14]=1;ram[107][15]=1;ram[107][16]=0;ram[107][17]=0;ram[107][18]=0;ram[107][19]=1;ram[107][20]=0;ram[107][21]=0;ram[107][22]=1;ram[107][23]=0;ram[107][24]=0;ram[107][25]=0;ram[107][26]=0;ram[107][27]=1;ram[107][28]=0;ram[107][29]=0;ram[107][30]=0;ram[107][31]=1;ram[107][32]=0;ram[107][33]=1;ram[107][34]=0;ram[107][35]=1;ram[107][36]=1;ram[107][37]=0;ram[107][38]=1;ram[107][39]=1;ram[107][40]=1;ram[107][41]=0;ram[107][42]=1;ram[107][43]=1;ram[107][44]=1;ram[107][45]=1;ram[107][46]=1;ram[107][47]=0;ram[107][48]=0;ram[107][49]=0;ram[107][50]=0;ram[107][51]=1;ram[107][52]=1;ram[107][53]=1;ram[107][54]=1;ram[107][55]=0;ram[107][56]=1;ram[107][57]=1;ram[107][58]=0;ram[107][59]=1;ram[107][60]=0;ram[107][61]=0;ram[107][62]=1;ram[107][63]=1;ram[107][64]=1;ram[107][65]=1;ram[107][66]=0;ram[107][67]=1;ram[107][68]=1;ram[107][69]=1;ram[107][70]=1;ram[107][71]=1;ram[107][72]=0;ram[107][73]=1;ram[107][74]=1;ram[107][75]=1;ram[107][76]=0;ram[107][77]=0;ram[107][78]=1;ram[107][79]=1;ram[107][80]=1;ram[107][81]=0;ram[107][82]=1;ram[107][83]=1;ram[107][84]=0;ram[107][85]=1;ram[107][86]=0;ram[107][87]=0;ram[107][88]=1;ram[107][89]=0;ram[107][90]=0;ram[107][91]=0;ram[107][92]=1;ram[107][93]=1;ram[107][94]=1;ram[107][95]=0;ram[107][96]=1;ram[107][97]=0;ram[107][98]=0;ram[107][99]=1;ram[107][100]=1;ram[107][101]=1;ram[107][102]=0;ram[107][103]=0;ram[107][104]=1;ram[107][105]=0;ram[107][106]=1;ram[107][107]=0;ram[107][108]=1;ram[107][109]=1;ram[107][110]=0;ram[107][111]=1;ram[107][112]=0;ram[107][113]=1;ram[107][114]=0;ram[107][115]=1;ram[107][116]=0;ram[107][117]=0;ram[107][118]=0;ram[107][119]=1;ram[107][120]=1;ram[107][121]=0;ram[107][122]=1;ram[107][123]=0;ram[107][124]=1;ram[107][125]=1;ram[107][126]=1;ram[107][127]=0;ram[107][128]=1;ram[107][129]=1;ram[107][130]=0;ram[107][131]=0;ram[107][132]=1;ram[107][133]=0;ram[107][134]=1;ram[107][135]=0;ram[107][136]=0;
        ram[108][0]=0;ram[108][1]=1;ram[108][2]=0;ram[108][3]=1;ram[108][4]=0;ram[108][5]=1;ram[108][6]=0;ram[108][7]=1;ram[108][8]=1;ram[108][9]=1;ram[108][10]=1;ram[108][11]=1;ram[108][12]=0;ram[108][13]=0;ram[108][14]=1;ram[108][15]=1;ram[108][16]=1;ram[108][17]=1;ram[108][18]=1;ram[108][19]=1;ram[108][20]=0;ram[108][21]=1;ram[108][22]=1;ram[108][23]=1;ram[108][24]=1;ram[108][25]=0;ram[108][26]=1;ram[108][27]=1;ram[108][28]=1;ram[108][29]=0;ram[108][30]=0;ram[108][31]=1;ram[108][32]=1;ram[108][33]=1;ram[108][34]=1;ram[108][35]=1;ram[108][36]=1;ram[108][37]=0;ram[108][38]=1;ram[108][39]=0;ram[108][40]=0;ram[108][41]=1;ram[108][42]=0;ram[108][43]=1;ram[108][44]=1;ram[108][45]=1;ram[108][46]=1;ram[108][47]=0;ram[108][48]=0;ram[108][49]=1;ram[108][50]=1;ram[108][51]=1;ram[108][52]=1;ram[108][53]=1;ram[108][54]=0;ram[108][55]=0;ram[108][56]=1;ram[108][57]=0;ram[108][58]=1;ram[108][59]=1;ram[108][60]=1;ram[108][61]=0;ram[108][62]=0;ram[108][63]=1;ram[108][64]=1;ram[108][65]=0;ram[108][66]=1;ram[108][67]=1;ram[108][68]=0;ram[108][69]=0;ram[108][70]=0;ram[108][71]=1;ram[108][72]=1;ram[108][73]=1;ram[108][74]=1;ram[108][75]=0;ram[108][76]=1;ram[108][77]=1;ram[108][78]=1;ram[108][79]=1;ram[108][80]=0;ram[108][81]=1;ram[108][82]=1;ram[108][83]=0;ram[108][84]=1;ram[108][85]=0;ram[108][86]=1;ram[108][87]=1;ram[108][88]=0;ram[108][89]=0;ram[108][90]=1;ram[108][91]=0;ram[108][92]=0;ram[108][93]=1;ram[108][94]=1;ram[108][95]=1;ram[108][96]=0;ram[108][97]=0;ram[108][98]=1;ram[108][99]=1;ram[108][100]=1;ram[108][101]=1;ram[108][102]=0;ram[108][103]=0;ram[108][104]=1;ram[108][105]=1;ram[108][106]=1;ram[108][107]=1;ram[108][108]=1;ram[108][109]=0;ram[108][110]=0;ram[108][111]=0;ram[108][112]=1;ram[108][113]=1;ram[108][114]=0;ram[108][115]=1;ram[108][116]=1;ram[108][117]=0;ram[108][118]=0;ram[108][119]=0;ram[108][120]=1;ram[108][121]=1;ram[108][122]=0;ram[108][123]=0;ram[108][124]=1;ram[108][125]=0;ram[108][126]=1;ram[108][127]=0;ram[108][128]=0;ram[108][129]=0;ram[108][130]=0;ram[108][131]=1;ram[108][132]=1;ram[108][133]=0;ram[108][134]=1;ram[108][135]=0;ram[108][136]=1;
        ram[109][0]=1;ram[109][1]=0;ram[109][2]=0;ram[109][3]=1;ram[109][4]=1;ram[109][5]=1;ram[109][6]=0;ram[109][7]=0;ram[109][8]=0;ram[109][9]=0;ram[109][10]=0;ram[109][11]=1;ram[109][12]=0;ram[109][13]=0;ram[109][14]=1;ram[109][15]=1;ram[109][16]=1;ram[109][17]=1;ram[109][18]=0;ram[109][19]=1;ram[109][20]=0;ram[109][21]=1;ram[109][22]=1;ram[109][23]=1;ram[109][24]=1;ram[109][25]=0;ram[109][26]=1;ram[109][27]=1;ram[109][28]=1;ram[109][29]=1;ram[109][30]=0;ram[109][31]=0;ram[109][32]=1;ram[109][33]=1;ram[109][34]=1;ram[109][35]=0;ram[109][36]=1;ram[109][37]=1;ram[109][38]=1;ram[109][39]=1;ram[109][40]=0;ram[109][41]=1;ram[109][42]=0;ram[109][43]=1;ram[109][44]=1;ram[109][45]=0;ram[109][46]=0;ram[109][47]=0;ram[109][48]=1;ram[109][49]=1;ram[109][50]=1;ram[109][51]=1;ram[109][52]=0;ram[109][53]=1;ram[109][54]=1;ram[109][55]=1;ram[109][56]=1;ram[109][57]=1;ram[109][58]=1;ram[109][59]=1;ram[109][60]=1;ram[109][61]=1;ram[109][62]=0;ram[109][63]=1;ram[109][64]=0;ram[109][65]=1;ram[109][66]=1;ram[109][67]=1;ram[109][68]=0;ram[109][69]=0;ram[109][70]=0;ram[109][71]=1;ram[109][72]=1;ram[109][73]=1;ram[109][74]=0;ram[109][75]=1;ram[109][76]=0;ram[109][77]=0;ram[109][78]=1;ram[109][79]=1;ram[109][80]=0;ram[109][81]=1;ram[109][82]=0;ram[109][83]=1;ram[109][84]=0;ram[109][85]=1;ram[109][86]=1;ram[109][87]=1;ram[109][88]=1;ram[109][89]=0;ram[109][90]=0;ram[109][91]=0;ram[109][92]=1;ram[109][93]=0;ram[109][94]=1;ram[109][95]=1;ram[109][96]=1;ram[109][97]=1;ram[109][98]=0;ram[109][99]=1;ram[109][100]=1;ram[109][101]=1;ram[109][102]=1;ram[109][103]=1;ram[109][104]=0;ram[109][105]=1;ram[109][106]=1;ram[109][107]=1;ram[109][108]=1;ram[109][109]=1;ram[109][110]=1;ram[109][111]=1;ram[109][112]=1;ram[109][113]=0;ram[109][114]=1;ram[109][115]=1;ram[109][116]=0;ram[109][117]=1;ram[109][118]=1;ram[109][119]=0;ram[109][120]=1;ram[109][121]=0;ram[109][122]=1;ram[109][123]=1;ram[109][124]=1;ram[109][125]=1;ram[109][126]=1;ram[109][127]=1;ram[109][128]=1;ram[109][129]=1;ram[109][130]=1;ram[109][131]=1;ram[109][132]=0;ram[109][133]=0;ram[109][134]=0;ram[109][135]=1;ram[109][136]=1;
        ram[110][0]=1;ram[110][1]=1;ram[110][2]=1;ram[110][3]=0;ram[110][4]=1;ram[110][5]=0;ram[110][6]=1;ram[110][7]=1;ram[110][8]=1;ram[110][9]=1;ram[110][10]=1;ram[110][11]=1;ram[110][12]=1;ram[110][13]=1;ram[110][14]=1;ram[110][15]=1;ram[110][16]=1;ram[110][17]=1;ram[110][18]=1;ram[110][19]=1;ram[110][20]=0;ram[110][21]=1;ram[110][22]=1;ram[110][23]=1;ram[110][24]=0;ram[110][25]=1;ram[110][26]=1;ram[110][27]=0;ram[110][28]=0;ram[110][29]=1;ram[110][30]=1;ram[110][31]=1;ram[110][32]=1;ram[110][33]=0;ram[110][34]=1;ram[110][35]=1;ram[110][36]=1;ram[110][37]=0;ram[110][38]=1;ram[110][39]=1;ram[110][40]=0;ram[110][41]=1;ram[110][42]=0;ram[110][43]=1;ram[110][44]=1;ram[110][45]=1;ram[110][46]=1;ram[110][47]=1;ram[110][48]=1;ram[110][49]=0;ram[110][50]=0;ram[110][51]=1;ram[110][52]=1;ram[110][53]=1;ram[110][54]=1;ram[110][55]=1;ram[110][56]=1;ram[110][57]=0;ram[110][58]=1;ram[110][59]=1;ram[110][60]=0;ram[110][61]=1;ram[110][62]=1;ram[110][63]=1;ram[110][64]=1;ram[110][65]=0;ram[110][66]=1;ram[110][67]=0;ram[110][68]=0;ram[110][69]=0;ram[110][70]=1;ram[110][71]=1;ram[110][72]=0;ram[110][73]=1;ram[110][74]=1;ram[110][75]=1;ram[110][76]=1;ram[110][77]=1;ram[110][78]=0;ram[110][79]=1;ram[110][80]=1;ram[110][81]=1;ram[110][82]=1;ram[110][83]=0;ram[110][84]=0;ram[110][85]=0;ram[110][86]=1;ram[110][87]=0;ram[110][88]=0;ram[110][89]=0;ram[110][90]=1;ram[110][91]=1;ram[110][92]=0;ram[110][93]=1;ram[110][94]=1;ram[110][95]=1;ram[110][96]=1;ram[110][97]=1;ram[110][98]=0;ram[110][99]=0;ram[110][100]=1;ram[110][101]=1;ram[110][102]=1;ram[110][103]=0;ram[110][104]=1;ram[110][105]=1;ram[110][106]=0;ram[110][107]=1;ram[110][108]=1;ram[110][109]=0;ram[110][110]=0;ram[110][111]=0;ram[110][112]=1;ram[110][113]=1;ram[110][114]=1;ram[110][115]=1;ram[110][116]=1;ram[110][117]=1;ram[110][118]=1;ram[110][119]=0;ram[110][120]=0;ram[110][121]=1;ram[110][122]=1;ram[110][123]=1;ram[110][124]=1;ram[110][125]=0;ram[110][126]=0;ram[110][127]=0;ram[110][128]=1;ram[110][129]=0;ram[110][130]=0;ram[110][131]=1;ram[110][132]=1;ram[110][133]=1;ram[110][134]=0;ram[110][135]=0;ram[110][136]=1;
        ram[111][0]=1;ram[111][1]=0;ram[111][2]=1;ram[111][3]=1;ram[111][4]=1;ram[111][5]=1;ram[111][6]=0;ram[111][7]=0;ram[111][8]=1;ram[111][9]=0;ram[111][10]=0;ram[111][11]=1;ram[111][12]=1;ram[111][13]=1;ram[111][14]=1;ram[111][15]=1;ram[111][16]=1;ram[111][17]=1;ram[111][18]=1;ram[111][19]=1;ram[111][20]=0;ram[111][21]=1;ram[111][22]=1;ram[111][23]=1;ram[111][24]=1;ram[111][25]=1;ram[111][26]=0;ram[111][27]=1;ram[111][28]=1;ram[111][29]=1;ram[111][30]=1;ram[111][31]=1;ram[111][32]=0;ram[111][33]=1;ram[111][34]=1;ram[111][35]=1;ram[111][36]=1;ram[111][37]=1;ram[111][38]=0;ram[111][39]=1;ram[111][40]=1;ram[111][41]=0;ram[111][42]=1;ram[111][43]=1;ram[111][44]=0;ram[111][45]=0;ram[111][46]=1;ram[111][47]=1;ram[111][48]=0;ram[111][49]=0;ram[111][50]=0;ram[111][51]=1;ram[111][52]=1;ram[111][53]=0;ram[111][54]=1;ram[111][55]=0;ram[111][56]=0;ram[111][57]=1;ram[111][58]=1;ram[111][59]=0;ram[111][60]=1;ram[111][61]=1;ram[111][62]=1;ram[111][63]=1;ram[111][64]=1;ram[111][65]=1;ram[111][66]=1;ram[111][67]=1;ram[111][68]=0;ram[111][69]=0;ram[111][70]=0;ram[111][71]=1;ram[111][72]=1;ram[111][73]=1;ram[111][74]=0;ram[111][75]=1;ram[111][76]=1;ram[111][77]=1;ram[111][78]=1;ram[111][79]=1;ram[111][80]=1;ram[111][81]=1;ram[111][82]=1;ram[111][83]=0;ram[111][84]=0;ram[111][85]=0;ram[111][86]=1;ram[111][87]=1;ram[111][88]=1;ram[111][89]=1;ram[111][90]=1;ram[111][91]=0;ram[111][92]=0;ram[111][93]=1;ram[111][94]=1;ram[111][95]=1;ram[111][96]=0;ram[111][97]=1;ram[111][98]=0;ram[111][99]=0;ram[111][100]=1;ram[111][101]=0;ram[111][102]=1;ram[111][103]=1;ram[111][104]=1;ram[111][105]=0;ram[111][106]=1;ram[111][107]=0;ram[111][108]=0;ram[111][109]=0;ram[111][110]=1;ram[111][111]=0;ram[111][112]=1;ram[111][113]=0;ram[111][114]=1;ram[111][115]=1;ram[111][116]=1;ram[111][117]=1;ram[111][118]=1;ram[111][119]=1;ram[111][120]=1;ram[111][121]=1;ram[111][122]=1;ram[111][123]=0;ram[111][124]=1;ram[111][125]=0;ram[111][126]=0;ram[111][127]=1;ram[111][128]=1;ram[111][129]=1;ram[111][130]=1;ram[111][131]=1;ram[111][132]=1;ram[111][133]=1;ram[111][134]=1;ram[111][135]=0;ram[111][136]=1;
        ram[112][0]=1;ram[112][1]=0;ram[112][2]=1;ram[112][3]=1;ram[112][4]=1;ram[112][5]=1;ram[112][6]=1;ram[112][7]=1;ram[112][8]=1;ram[112][9]=1;ram[112][10]=0;ram[112][11]=0;ram[112][12]=1;ram[112][13]=1;ram[112][14]=1;ram[112][15]=1;ram[112][16]=0;ram[112][17]=1;ram[112][18]=1;ram[112][19]=1;ram[112][20]=1;ram[112][21]=1;ram[112][22]=1;ram[112][23]=0;ram[112][24]=0;ram[112][25]=1;ram[112][26]=1;ram[112][27]=1;ram[112][28]=0;ram[112][29]=1;ram[112][30]=1;ram[112][31]=1;ram[112][32]=0;ram[112][33]=1;ram[112][34]=1;ram[112][35]=0;ram[112][36]=0;ram[112][37]=1;ram[112][38]=1;ram[112][39]=0;ram[112][40]=1;ram[112][41]=1;ram[112][42]=1;ram[112][43]=1;ram[112][44]=1;ram[112][45]=1;ram[112][46]=1;ram[112][47]=1;ram[112][48]=1;ram[112][49]=0;ram[112][50]=1;ram[112][51]=0;ram[112][52]=1;ram[112][53]=1;ram[112][54]=0;ram[112][55]=0;ram[112][56]=0;ram[112][57]=1;ram[112][58]=1;ram[112][59]=0;ram[112][60]=0;ram[112][61]=1;ram[112][62]=1;ram[112][63]=0;ram[112][64]=1;ram[112][65]=1;ram[112][66]=1;ram[112][67]=1;ram[112][68]=0;ram[112][69]=1;ram[112][70]=1;ram[112][71]=1;ram[112][72]=1;ram[112][73]=1;ram[112][74]=1;ram[112][75]=1;ram[112][76]=1;ram[112][77]=1;ram[112][78]=1;ram[112][79]=1;ram[112][80]=1;ram[112][81]=0;ram[112][82]=1;ram[112][83]=1;ram[112][84]=1;ram[112][85]=1;ram[112][86]=1;ram[112][87]=0;ram[112][88]=1;ram[112][89]=1;ram[112][90]=0;ram[112][91]=1;ram[112][92]=0;ram[112][93]=1;ram[112][94]=1;ram[112][95]=1;ram[112][96]=0;ram[112][97]=1;ram[112][98]=0;ram[112][99]=1;ram[112][100]=1;ram[112][101]=0;ram[112][102]=0;ram[112][103]=1;ram[112][104]=1;ram[112][105]=1;ram[112][106]=1;ram[112][107]=1;ram[112][108]=1;ram[112][109]=1;ram[112][110]=1;ram[112][111]=0;ram[112][112]=1;ram[112][113]=1;ram[112][114]=0;ram[112][115]=0;ram[112][116]=1;ram[112][117]=1;ram[112][118]=1;ram[112][119]=1;ram[112][120]=1;ram[112][121]=1;ram[112][122]=1;ram[112][123]=1;ram[112][124]=0;ram[112][125]=0;ram[112][126]=1;ram[112][127]=0;ram[112][128]=0;ram[112][129]=1;ram[112][130]=1;ram[112][131]=1;ram[112][132]=1;ram[112][133]=1;ram[112][134]=1;ram[112][135]=0;ram[112][136]=0;
        ram[113][0]=1;ram[113][1]=0;ram[113][2]=1;ram[113][3]=0;ram[113][4]=1;ram[113][5]=1;ram[113][6]=0;ram[113][7]=1;ram[113][8]=1;ram[113][9]=1;ram[113][10]=1;ram[113][11]=1;ram[113][12]=0;ram[113][13]=0;ram[113][14]=0;ram[113][15]=1;ram[113][16]=1;ram[113][17]=1;ram[113][18]=0;ram[113][19]=1;ram[113][20]=0;ram[113][21]=0;ram[113][22]=1;ram[113][23]=1;ram[113][24]=1;ram[113][25]=1;ram[113][26]=0;ram[113][27]=0;ram[113][28]=1;ram[113][29]=0;ram[113][30]=0;ram[113][31]=0;ram[113][32]=1;ram[113][33]=0;ram[113][34]=0;ram[113][35]=1;ram[113][36]=1;ram[113][37]=1;ram[113][38]=1;ram[113][39]=0;ram[113][40]=0;ram[113][41]=1;ram[113][42]=0;ram[113][43]=1;ram[113][44]=0;ram[113][45]=1;ram[113][46]=1;ram[113][47]=1;ram[113][48]=0;ram[113][49]=1;ram[113][50]=1;ram[113][51]=1;ram[113][52]=1;ram[113][53]=1;ram[113][54]=1;ram[113][55]=0;ram[113][56]=1;ram[113][57]=0;ram[113][58]=0;ram[113][59]=1;ram[113][60]=1;ram[113][61]=0;ram[113][62]=1;ram[113][63]=1;ram[113][64]=1;ram[113][65]=0;ram[113][66]=1;ram[113][67]=0;ram[113][68]=1;ram[113][69]=0;ram[113][70]=0;ram[113][71]=0;ram[113][72]=1;ram[113][73]=0;ram[113][74]=1;ram[113][75]=1;ram[113][76]=1;ram[113][77]=0;ram[113][78]=1;ram[113][79]=1;ram[113][80]=1;ram[113][81]=1;ram[113][82]=0;ram[113][83]=1;ram[113][84]=1;ram[113][85]=1;ram[113][86]=0;ram[113][87]=1;ram[113][88]=1;ram[113][89]=0;ram[113][90]=1;ram[113][91]=0;ram[113][92]=1;ram[113][93]=1;ram[113][94]=1;ram[113][95]=1;ram[113][96]=1;ram[113][97]=1;ram[113][98]=1;ram[113][99]=1;ram[113][100]=1;ram[113][101]=1;ram[113][102]=0;ram[113][103]=1;ram[113][104]=1;ram[113][105]=0;ram[113][106]=1;ram[113][107]=0;ram[113][108]=1;ram[113][109]=1;ram[113][110]=1;ram[113][111]=1;ram[113][112]=1;ram[113][113]=1;ram[113][114]=1;ram[113][115]=1;ram[113][116]=1;ram[113][117]=0;ram[113][118]=0;ram[113][119]=0;ram[113][120]=1;ram[113][121]=0;ram[113][122]=1;ram[113][123]=1;ram[113][124]=0;ram[113][125]=1;ram[113][126]=1;ram[113][127]=0;ram[113][128]=1;ram[113][129]=0;ram[113][130]=0;ram[113][131]=0;ram[113][132]=1;ram[113][133]=1;ram[113][134]=1;ram[113][135]=1;ram[113][136]=1;
        ram[114][0]=0;ram[114][1]=0;ram[114][2]=1;ram[114][3]=1;ram[114][4]=1;ram[114][5]=0;ram[114][6]=0;ram[114][7]=1;ram[114][8]=1;ram[114][9]=1;ram[114][10]=0;ram[114][11]=1;ram[114][12]=0;ram[114][13]=1;ram[114][14]=1;ram[114][15]=1;ram[114][16]=1;ram[114][17]=0;ram[114][18]=1;ram[114][19]=1;ram[114][20]=1;ram[114][21]=0;ram[114][22]=1;ram[114][23]=1;ram[114][24]=0;ram[114][25]=0;ram[114][26]=1;ram[114][27]=1;ram[114][28]=0;ram[114][29]=1;ram[114][30]=0;ram[114][31]=1;ram[114][32]=0;ram[114][33]=1;ram[114][34]=0;ram[114][35]=1;ram[114][36]=1;ram[114][37]=1;ram[114][38]=0;ram[114][39]=1;ram[114][40]=0;ram[114][41]=1;ram[114][42]=1;ram[114][43]=1;ram[114][44]=1;ram[114][45]=1;ram[114][46]=1;ram[114][47]=1;ram[114][48]=1;ram[114][49]=1;ram[114][50]=0;ram[114][51]=0;ram[114][52]=1;ram[114][53]=0;ram[114][54]=1;ram[114][55]=0;ram[114][56]=0;ram[114][57]=1;ram[114][58]=0;ram[114][59]=1;ram[114][60]=1;ram[114][61]=1;ram[114][62]=0;ram[114][63]=0;ram[114][64]=1;ram[114][65]=1;ram[114][66]=0;ram[114][67]=0;ram[114][68]=0;ram[114][69]=1;ram[114][70]=1;ram[114][71]=0;ram[114][72]=0;ram[114][73]=1;ram[114][74]=0;ram[114][75]=1;ram[114][76]=0;ram[114][77]=0;ram[114][78]=1;ram[114][79]=0;ram[114][80]=0;ram[114][81]=0;ram[114][82]=1;ram[114][83]=1;ram[114][84]=1;ram[114][85]=1;ram[114][86]=0;ram[114][87]=0;ram[114][88]=1;ram[114][89]=0;ram[114][90]=1;ram[114][91]=1;ram[114][92]=0;ram[114][93]=1;ram[114][94]=1;ram[114][95]=0;ram[114][96]=1;ram[114][97]=1;ram[114][98]=1;ram[114][99]=1;ram[114][100]=1;ram[114][101]=1;ram[114][102]=0;ram[114][103]=0;ram[114][104]=1;ram[114][105]=0;ram[114][106]=0;ram[114][107]=1;ram[114][108]=1;ram[114][109]=1;ram[114][110]=0;ram[114][111]=0;ram[114][112]=0;ram[114][113]=1;ram[114][114]=1;ram[114][115]=1;ram[114][116]=0;ram[114][117]=1;ram[114][118]=0;ram[114][119]=1;ram[114][120]=1;ram[114][121]=1;ram[114][122]=0;ram[114][123]=1;ram[114][124]=0;ram[114][125]=1;ram[114][126]=1;ram[114][127]=1;ram[114][128]=0;ram[114][129]=0;ram[114][130]=0;ram[114][131]=1;ram[114][132]=1;ram[114][133]=1;ram[114][134]=1;ram[114][135]=1;ram[114][136]=0;
        ram[115][0]=0;ram[115][1]=1;ram[115][2]=0;ram[115][3]=1;ram[115][4]=1;ram[115][5]=0;ram[115][6]=1;ram[115][7]=1;ram[115][8]=1;ram[115][9]=1;ram[115][10]=0;ram[115][11]=1;ram[115][12]=1;ram[115][13]=1;ram[115][14]=1;ram[115][15]=0;ram[115][16]=0;ram[115][17]=1;ram[115][18]=1;ram[115][19]=1;ram[115][20]=0;ram[115][21]=1;ram[115][22]=0;ram[115][23]=1;ram[115][24]=1;ram[115][25]=1;ram[115][26]=1;ram[115][27]=1;ram[115][28]=1;ram[115][29]=0;ram[115][30]=1;ram[115][31]=0;ram[115][32]=0;ram[115][33]=1;ram[115][34]=1;ram[115][35]=1;ram[115][36]=0;ram[115][37]=1;ram[115][38]=1;ram[115][39]=0;ram[115][40]=1;ram[115][41]=1;ram[115][42]=1;ram[115][43]=1;ram[115][44]=1;ram[115][45]=1;ram[115][46]=1;ram[115][47]=1;ram[115][48]=0;ram[115][49]=0;ram[115][50]=1;ram[115][51]=1;ram[115][52]=1;ram[115][53]=0;ram[115][54]=0;ram[115][55]=1;ram[115][56]=0;ram[115][57]=0;ram[115][58]=1;ram[115][59]=1;ram[115][60]=1;ram[115][61]=0;ram[115][62]=0;ram[115][63]=0;ram[115][64]=1;ram[115][65]=1;ram[115][66]=1;ram[115][67]=0;ram[115][68]=1;ram[115][69]=1;ram[115][70]=0;ram[115][71]=1;ram[115][72]=1;ram[115][73]=1;ram[115][74]=0;ram[115][75]=0;ram[115][76]=0;ram[115][77]=0;ram[115][78]=1;ram[115][79]=1;ram[115][80]=1;ram[115][81]=1;ram[115][82]=1;ram[115][83]=1;ram[115][84]=1;ram[115][85]=1;ram[115][86]=1;ram[115][87]=1;ram[115][88]=1;ram[115][89]=1;ram[115][90]=1;ram[115][91]=0;ram[115][92]=0;ram[115][93]=1;ram[115][94]=1;ram[115][95]=0;ram[115][96]=1;ram[115][97]=1;ram[115][98]=1;ram[115][99]=1;ram[115][100]=0;ram[115][101]=0;ram[115][102]=1;ram[115][103]=1;ram[115][104]=1;ram[115][105]=1;ram[115][106]=0;ram[115][107]=1;ram[115][108]=0;ram[115][109]=0;ram[115][110]=1;ram[115][111]=1;ram[115][112]=1;ram[115][113]=1;ram[115][114]=0;ram[115][115]=1;ram[115][116]=0;ram[115][117]=1;ram[115][118]=0;ram[115][119]=0;ram[115][120]=1;ram[115][121]=1;ram[115][122]=1;ram[115][123]=1;ram[115][124]=1;ram[115][125]=1;ram[115][126]=1;ram[115][127]=1;ram[115][128]=0;ram[115][129]=1;ram[115][130]=0;ram[115][131]=1;ram[115][132]=0;ram[115][133]=1;ram[115][134]=0;ram[115][135]=1;ram[115][136]=1;
        ram[116][0]=1;ram[116][1]=1;ram[116][2]=1;ram[116][3]=1;ram[116][4]=0;ram[116][5]=1;ram[116][6]=1;ram[116][7]=1;ram[116][8]=1;ram[116][9]=0;ram[116][10]=1;ram[116][11]=0;ram[116][12]=0;ram[116][13]=1;ram[116][14]=1;ram[116][15]=1;ram[116][16]=0;ram[116][17]=0;ram[116][18]=1;ram[116][19]=1;ram[116][20]=1;ram[116][21]=1;ram[116][22]=0;ram[116][23]=1;ram[116][24]=1;ram[116][25]=0;ram[116][26]=1;ram[116][27]=1;ram[116][28]=0;ram[116][29]=1;ram[116][30]=0;ram[116][31]=0;ram[116][32]=1;ram[116][33]=1;ram[116][34]=1;ram[116][35]=1;ram[116][36]=1;ram[116][37]=1;ram[116][38]=0;ram[116][39]=0;ram[116][40]=0;ram[116][41]=0;ram[116][42]=1;ram[116][43]=1;ram[116][44]=1;ram[116][45]=1;ram[116][46]=1;ram[116][47]=0;ram[116][48]=0;ram[116][49]=1;ram[116][50]=1;ram[116][51]=1;ram[116][52]=1;ram[116][53]=0;ram[116][54]=0;ram[116][55]=1;ram[116][56]=1;ram[116][57]=0;ram[116][58]=1;ram[116][59]=1;ram[116][60]=1;ram[116][61]=1;ram[116][62]=1;ram[116][63]=1;ram[116][64]=0;ram[116][65]=1;ram[116][66]=0;ram[116][67]=0;ram[116][68]=0;ram[116][69]=1;ram[116][70]=0;ram[116][71]=1;ram[116][72]=1;ram[116][73]=0;ram[116][74]=0;ram[116][75]=1;ram[116][76]=1;ram[116][77]=0;ram[116][78]=1;ram[116][79]=1;ram[116][80]=1;ram[116][81]=1;ram[116][82]=1;ram[116][83]=1;ram[116][84]=1;ram[116][85]=1;ram[116][86]=0;ram[116][87]=1;ram[116][88]=0;ram[116][89]=1;ram[116][90]=1;ram[116][91]=1;ram[116][92]=1;ram[116][93]=1;ram[116][94]=0;ram[116][95]=0;ram[116][96]=0;ram[116][97]=0;ram[116][98]=0;ram[116][99]=1;ram[116][100]=0;ram[116][101]=0;ram[116][102]=1;ram[116][103]=0;ram[116][104]=1;ram[116][105]=1;ram[116][106]=1;ram[116][107]=1;ram[116][108]=0;ram[116][109]=1;ram[116][110]=1;ram[116][111]=1;ram[116][112]=0;ram[116][113]=1;ram[116][114]=1;ram[116][115]=1;ram[116][116]=0;ram[116][117]=1;ram[116][118]=1;ram[116][119]=0;ram[116][120]=0;ram[116][121]=1;ram[116][122]=1;ram[116][123]=1;ram[116][124]=1;ram[116][125]=1;ram[116][126]=1;ram[116][127]=1;ram[116][128]=1;ram[116][129]=1;ram[116][130]=0;ram[116][131]=1;ram[116][132]=0;ram[116][133]=0;ram[116][134]=1;ram[116][135]=1;ram[116][136]=0;
        ram[117][0]=0;ram[117][1]=0;ram[117][2]=1;ram[117][3]=1;ram[117][4]=1;ram[117][5]=1;ram[117][6]=1;ram[117][7]=1;ram[117][8]=1;ram[117][9]=1;ram[117][10]=0;ram[117][11]=1;ram[117][12]=1;ram[117][13]=0;ram[117][14]=0;ram[117][15]=1;ram[117][16]=1;ram[117][17]=1;ram[117][18]=0;ram[117][19]=1;ram[117][20]=1;ram[117][21]=0;ram[117][22]=1;ram[117][23]=0;ram[117][24]=0;ram[117][25]=0;ram[117][26]=1;ram[117][27]=1;ram[117][28]=1;ram[117][29]=0;ram[117][30]=0;ram[117][31]=1;ram[117][32]=0;ram[117][33]=0;ram[117][34]=1;ram[117][35]=0;ram[117][36]=0;ram[117][37]=1;ram[117][38]=1;ram[117][39]=1;ram[117][40]=0;ram[117][41]=0;ram[117][42]=1;ram[117][43]=1;ram[117][44]=1;ram[117][45]=1;ram[117][46]=1;ram[117][47]=0;ram[117][48]=1;ram[117][49]=1;ram[117][50]=1;ram[117][51]=0;ram[117][52]=0;ram[117][53]=1;ram[117][54]=1;ram[117][55]=1;ram[117][56]=1;ram[117][57]=0;ram[117][58]=1;ram[117][59]=0;ram[117][60]=1;ram[117][61]=0;ram[117][62]=1;ram[117][63]=0;ram[117][64]=1;ram[117][65]=0;ram[117][66]=1;ram[117][67]=1;ram[117][68]=0;ram[117][69]=1;ram[117][70]=1;ram[117][71]=1;ram[117][72]=1;ram[117][73]=1;ram[117][74]=1;ram[117][75]=0;ram[117][76]=1;ram[117][77]=1;ram[117][78]=0;ram[117][79]=1;ram[117][80]=1;ram[117][81]=0;ram[117][82]=1;ram[117][83]=1;ram[117][84]=1;ram[117][85]=1;ram[117][86]=0;ram[117][87]=1;ram[117][88]=1;ram[117][89]=0;ram[117][90]=0;ram[117][91]=0;ram[117][92]=1;ram[117][93]=0;ram[117][94]=1;ram[117][95]=1;ram[117][96]=1;ram[117][97]=1;ram[117][98]=1;ram[117][99]=1;ram[117][100]=0;ram[117][101]=1;ram[117][102]=0;ram[117][103]=1;ram[117][104]=0;ram[117][105]=1;ram[117][106]=1;ram[117][107]=1;ram[117][108]=0;ram[117][109]=0;ram[117][110]=0;ram[117][111]=1;ram[117][112]=1;ram[117][113]=1;ram[117][114]=1;ram[117][115]=0;ram[117][116]=1;ram[117][117]=1;ram[117][118]=1;ram[117][119]=0;ram[117][120]=1;ram[117][121]=1;ram[117][122]=1;ram[117][123]=0;ram[117][124]=1;ram[117][125]=0;ram[117][126]=1;ram[117][127]=1;ram[117][128]=0;ram[117][129]=0;ram[117][130]=1;ram[117][131]=1;ram[117][132]=1;ram[117][133]=1;ram[117][134]=0;ram[117][135]=0;ram[117][136]=1;
        ram[118][0]=0;ram[118][1]=0;ram[118][2]=1;ram[118][3]=1;ram[118][4]=0;ram[118][5]=1;ram[118][6]=0;ram[118][7]=0;ram[118][8]=1;ram[118][9]=1;ram[118][10]=1;ram[118][11]=1;ram[118][12]=1;ram[118][13]=1;ram[118][14]=1;ram[118][15]=1;ram[118][16]=1;ram[118][17]=1;ram[118][18]=1;ram[118][19]=1;ram[118][20]=1;ram[118][21]=1;ram[118][22]=0;ram[118][23]=1;ram[118][24]=1;ram[118][25]=1;ram[118][26]=1;ram[118][27]=0;ram[118][28]=1;ram[118][29]=1;ram[118][30]=1;ram[118][31]=0;ram[118][32]=1;ram[118][33]=1;ram[118][34]=1;ram[118][35]=1;ram[118][36]=1;ram[118][37]=1;ram[118][38]=0;ram[118][39]=1;ram[118][40]=1;ram[118][41]=1;ram[118][42]=1;ram[118][43]=1;ram[118][44]=0;ram[118][45]=0;ram[118][46]=1;ram[118][47]=1;ram[118][48]=0;ram[118][49]=0;ram[118][50]=0;ram[118][51]=1;ram[118][52]=1;ram[118][53]=0;ram[118][54]=0;ram[118][55]=0;ram[118][56]=1;ram[118][57]=1;ram[118][58]=1;ram[118][59]=0;ram[118][60]=1;ram[118][61]=0;ram[118][62]=0;ram[118][63]=1;ram[118][64]=1;ram[118][65]=0;ram[118][66]=1;ram[118][67]=0;ram[118][68]=1;ram[118][69]=1;ram[118][70]=0;ram[118][71]=1;ram[118][72]=0;ram[118][73]=0;ram[118][74]=0;ram[118][75]=1;ram[118][76]=0;ram[118][77]=1;ram[118][78]=1;ram[118][79]=0;ram[118][80]=1;ram[118][81]=1;ram[118][82]=0;ram[118][83]=0;ram[118][84]=1;ram[118][85]=1;ram[118][86]=1;ram[118][87]=1;ram[118][88]=0;ram[118][89]=1;ram[118][90]=0;ram[118][91]=0;ram[118][92]=1;ram[118][93]=1;ram[118][94]=1;ram[118][95]=0;ram[118][96]=0;ram[118][97]=0;ram[118][98]=0;ram[118][99]=1;ram[118][100]=0;ram[118][101]=1;ram[118][102]=1;ram[118][103]=1;ram[118][104]=1;ram[118][105]=0;ram[118][106]=1;ram[118][107]=0;ram[118][108]=0;ram[118][109]=0;ram[118][110]=1;ram[118][111]=1;ram[118][112]=1;ram[118][113]=1;ram[118][114]=0;ram[118][115]=1;ram[118][116]=1;ram[118][117]=1;ram[118][118]=0;ram[118][119]=0;ram[118][120]=1;ram[118][121]=1;ram[118][122]=0;ram[118][123]=0;ram[118][124]=1;ram[118][125]=1;ram[118][126]=1;ram[118][127]=1;ram[118][128]=1;ram[118][129]=0;ram[118][130]=1;ram[118][131]=1;ram[118][132]=1;ram[118][133]=1;ram[118][134]=1;ram[118][135]=1;ram[118][136]=1;
        ram[119][0]=1;ram[119][1]=1;ram[119][2]=1;ram[119][3]=1;ram[119][4]=1;ram[119][5]=0;ram[119][6]=1;ram[119][7]=1;ram[119][8]=1;ram[119][9]=0;ram[119][10]=0;ram[119][11]=1;ram[119][12]=1;ram[119][13]=0;ram[119][14]=0;ram[119][15]=1;ram[119][16]=0;ram[119][17]=1;ram[119][18]=0;ram[119][19]=0;ram[119][20]=0;ram[119][21]=1;ram[119][22]=0;ram[119][23]=0;ram[119][24]=1;ram[119][25]=1;ram[119][26]=0;ram[119][27]=0;ram[119][28]=0;ram[119][29]=0;ram[119][30]=0;ram[119][31]=1;ram[119][32]=0;ram[119][33]=1;ram[119][34]=0;ram[119][35]=1;ram[119][36]=1;ram[119][37]=0;ram[119][38]=0;ram[119][39]=0;ram[119][40]=1;ram[119][41]=0;ram[119][42]=1;ram[119][43]=0;ram[119][44]=1;ram[119][45]=0;ram[119][46]=1;ram[119][47]=1;ram[119][48]=0;ram[119][49]=1;ram[119][50]=0;ram[119][51]=1;ram[119][52]=1;ram[119][53]=0;ram[119][54]=0;ram[119][55]=1;ram[119][56]=1;ram[119][57]=1;ram[119][58]=1;ram[119][59]=0;ram[119][60]=0;ram[119][61]=1;ram[119][62]=1;ram[119][63]=1;ram[119][64]=1;ram[119][65]=1;ram[119][66]=1;ram[119][67]=1;ram[119][68]=1;ram[119][69]=0;ram[119][70]=1;ram[119][71]=0;ram[119][72]=1;ram[119][73]=1;ram[119][74]=1;ram[119][75]=1;ram[119][76]=1;ram[119][77]=1;ram[119][78]=0;ram[119][79]=1;ram[119][80]=1;ram[119][81]=1;ram[119][82]=0;ram[119][83]=1;ram[119][84]=1;ram[119][85]=1;ram[119][86]=1;ram[119][87]=1;ram[119][88]=0;ram[119][89]=0;ram[119][90]=0;ram[119][91]=1;ram[119][92]=1;ram[119][93]=0;ram[119][94]=1;ram[119][95]=0;ram[119][96]=1;ram[119][97]=1;ram[119][98]=1;ram[119][99]=0;ram[119][100]=0;ram[119][101]=1;ram[119][102]=1;ram[119][103]=1;ram[119][104]=1;ram[119][105]=0;ram[119][106]=1;ram[119][107]=1;ram[119][108]=1;ram[119][109]=0;ram[119][110]=1;ram[119][111]=1;ram[119][112]=0;ram[119][113]=1;ram[119][114]=1;ram[119][115]=0;ram[119][116]=1;ram[119][117]=1;ram[119][118]=0;ram[119][119]=1;ram[119][120]=1;ram[119][121]=0;ram[119][122]=1;ram[119][123]=1;ram[119][124]=1;ram[119][125]=1;ram[119][126]=1;ram[119][127]=1;ram[119][128]=0;ram[119][129]=0;ram[119][130]=1;ram[119][131]=1;ram[119][132]=0;ram[119][133]=1;ram[119][134]=0;ram[119][135]=1;ram[119][136]=1;
        ram[120][0]=1;ram[120][1]=1;ram[120][2]=1;ram[120][3]=1;ram[120][4]=1;ram[120][5]=1;ram[120][6]=1;ram[120][7]=1;ram[120][8]=0;ram[120][9]=0;ram[120][10]=1;ram[120][11]=1;ram[120][12]=1;ram[120][13]=1;ram[120][14]=1;ram[120][15]=1;ram[120][16]=0;ram[120][17]=1;ram[120][18]=0;ram[120][19]=0;ram[120][20]=1;ram[120][21]=0;ram[120][22]=1;ram[120][23]=0;ram[120][24]=1;ram[120][25]=0;ram[120][26]=1;ram[120][27]=1;ram[120][28]=1;ram[120][29]=1;ram[120][30]=1;ram[120][31]=1;ram[120][32]=1;ram[120][33]=0;ram[120][34]=0;ram[120][35]=1;ram[120][36]=0;ram[120][37]=1;ram[120][38]=1;ram[120][39]=1;ram[120][40]=1;ram[120][41]=1;ram[120][42]=0;ram[120][43]=1;ram[120][44]=0;ram[120][45]=0;ram[120][46]=1;ram[120][47]=1;ram[120][48]=1;ram[120][49]=0;ram[120][50]=1;ram[120][51]=1;ram[120][52]=1;ram[120][53]=1;ram[120][54]=1;ram[120][55]=1;ram[120][56]=1;ram[120][57]=1;ram[120][58]=1;ram[120][59]=1;ram[120][60]=1;ram[120][61]=1;ram[120][62]=1;ram[120][63]=0;ram[120][64]=1;ram[120][65]=1;ram[120][66]=0;ram[120][67]=0;ram[120][68]=1;ram[120][69]=0;ram[120][70]=0;ram[120][71]=1;ram[120][72]=0;ram[120][73]=1;ram[120][74]=1;ram[120][75]=1;ram[120][76]=1;ram[120][77]=1;ram[120][78]=1;ram[120][79]=1;ram[120][80]=0;ram[120][81]=1;ram[120][82]=0;ram[120][83]=1;ram[120][84]=0;ram[120][85]=1;ram[120][86]=0;ram[120][87]=1;ram[120][88]=1;ram[120][89]=1;ram[120][90]=0;ram[120][91]=1;ram[120][92]=0;ram[120][93]=0;ram[120][94]=1;ram[120][95]=1;ram[120][96]=1;ram[120][97]=1;ram[120][98]=1;ram[120][99]=1;ram[120][100]=1;ram[120][101]=0;ram[120][102]=0;ram[120][103]=1;ram[120][104]=1;ram[120][105]=1;ram[120][106]=1;ram[120][107]=0;ram[120][108]=0;ram[120][109]=1;ram[120][110]=1;ram[120][111]=1;ram[120][112]=1;ram[120][113]=1;ram[120][114]=0;ram[120][115]=1;ram[120][116]=1;ram[120][117]=1;ram[120][118]=0;ram[120][119]=1;ram[120][120]=1;ram[120][121]=1;ram[120][122]=0;ram[120][123]=1;ram[120][124]=1;ram[120][125]=1;ram[120][126]=1;ram[120][127]=1;ram[120][128]=1;ram[120][129]=1;ram[120][130]=1;ram[120][131]=1;ram[120][132]=0;ram[120][133]=0;ram[120][134]=0;ram[120][135]=1;ram[120][136]=1;
        ram[121][0]=0;ram[121][1]=0;ram[121][2]=1;ram[121][3]=1;ram[121][4]=0;ram[121][5]=1;ram[121][6]=1;ram[121][7]=0;ram[121][8]=0;ram[121][9]=1;ram[121][10]=1;ram[121][11]=1;ram[121][12]=0;ram[121][13]=1;ram[121][14]=1;ram[121][15]=1;ram[121][16]=1;ram[121][17]=1;ram[121][18]=1;ram[121][19]=1;ram[121][20]=0;ram[121][21]=1;ram[121][22]=1;ram[121][23]=0;ram[121][24]=1;ram[121][25]=1;ram[121][26]=1;ram[121][27]=1;ram[121][28]=1;ram[121][29]=0;ram[121][30]=1;ram[121][31]=0;ram[121][32]=1;ram[121][33]=1;ram[121][34]=0;ram[121][35]=0;ram[121][36]=1;ram[121][37]=0;ram[121][38]=1;ram[121][39]=1;ram[121][40]=1;ram[121][41]=1;ram[121][42]=1;ram[121][43]=1;ram[121][44]=1;ram[121][45]=0;ram[121][46]=1;ram[121][47]=0;ram[121][48]=0;ram[121][49]=1;ram[121][50]=1;ram[121][51]=1;ram[121][52]=1;ram[121][53]=1;ram[121][54]=0;ram[121][55]=0;ram[121][56]=0;ram[121][57]=1;ram[121][58]=1;ram[121][59]=1;ram[121][60]=1;ram[121][61]=1;ram[121][62]=0;ram[121][63]=0;ram[121][64]=0;ram[121][65]=1;ram[121][66]=1;ram[121][67]=1;ram[121][68]=1;ram[121][69]=1;ram[121][70]=1;ram[121][71]=1;ram[121][72]=0;ram[121][73]=0;ram[121][74]=1;ram[121][75]=1;ram[121][76]=1;ram[121][77]=1;ram[121][78]=1;ram[121][79]=1;ram[121][80]=1;ram[121][81]=1;ram[121][82]=1;ram[121][83]=0;ram[121][84]=1;ram[121][85]=1;ram[121][86]=1;ram[121][87]=1;ram[121][88]=0;ram[121][89]=1;ram[121][90]=1;ram[121][91]=1;ram[121][92]=1;ram[121][93]=1;ram[121][94]=1;ram[121][95]=0;ram[121][96]=1;ram[121][97]=1;ram[121][98]=0;ram[121][99]=0;ram[121][100]=1;ram[121][101]=0;ram[121][102]=1;ram[121][103]=1;ram[121][104]=1;ram[121][105]=1;ram[121][106]=1;ram[121][107]=1;ram[121][108]=1;ram[121][109]=1;ram[121][110]=1;ram[121][111]=1;ram[121][112]=1;ram[121][113]=1;ram[121][114]=1;ram[121][115]=1;ram[121][116]=1;ram[121][117]=0;ram[121][118]=1;ram[121][119]=1;ram[121][120]=1;ram[121][121]=0;ram[121][122]=1;ram[121][123]=1;ram[121][124]=0;ram[121][125]=1;ram[121][126]=0;ram[121][127]=0;ram[121][128]=1;ram[121][129]=1;ram[121][130]=1;ram[121][131]=1;ram[121][132]=1;ram[121][133]=1;ram[121][134]=1;ram[121][135]=1;ram[121][136]=1;
        ram[122][0]=0;ram[122][1]=0;ram[122][2]=1;ram[122][3]=1;ram[122][4]=1;ram[122][5]=1;ram[122][6]=0;ram[122][7]=1;ram[122][8]=1;ram[122][9]=1;ram[122][10]=1;ram[122][11]=0;ram[122][12]=1;ram[122][13]=1;ram[122][14]=1;ram[122][15]=0;ram[122][16]=0;ram[122][17]=1;ram[122][18]=1;ram[122][19]=1;ram[122][20]=0;ram[122][21]=1;ram[122][22]=1;ram[122][23]=0;ram[122][24]=0;ram[122][25]=1;ram[122][26]=1;ram[122][27]=1;ram[122][28]=1;ram[122][29]=1;ram[122][30]=1;ram[122][31]=0;ram[122][32]=1;ram[122][33]=1;ram[122][34]=0;ram[122][35]=1;ram[122][36]=0;ram[122][37]=0;ram[122][38]=0;ram[122][39]=1;ram[122][40]=0;ram[122][41]=0;ram[122][42]=1;ram[122][43]=1;ram[122][44]=1;ram[122][45]=1;ram[122][46]=0;ram[122][47]=1;ram[122][48]=0;ram[122][49]=1;ram[122][50]=1;ram[122][51]=1;ram[122][52]=0;ram[122][53]=1;ram[122][54]=1;ram[122][55]=1;ram[122][56]=1;ram[122][57]=1;ram[122][58]=0;ram[122][59]=1;ram[122][60]=1;ram[122][61]=0;ram[122][62]=0;ram[122][63]=1;ram[122][64]=1;ram[122][65]=1;ram[122][66]=0;ram[122][67]=1;ram[122][68]=1;ram[122][69]=0;ram[122][70]=0;ram[122][71]=1;ram[122][72]=1;ram[122][73]=1;ram[122][74]=1;ram[122][75]=0;ram[122][76]=1;ram[122][77]=0;ram[122][78]=0;ram[122][79]=0;ram[122][80]=1;ram[122][81]=1;ram[122][82]=1;ram[122][83]=0;ram[122][84]=1;ram[122][85]=1;ram[122][86]=1;ram[122][87]=0;ram[122][88]=1;ram[122][89]=1;ram[122][90]=1;ram[122][91]=1;ram[122][92]=1;ram[122][93]=1;ram[122][94]=1;ram[122][95]=1;ram[122][96]=1;ram[122][97]=1;ram[122][98]=1;ram[122][99]=0;ram[122][100]=1;ram[122][101]=1;ram[122][102]=1;ram[122][103]=0;ram[122][104]=0;ram[122][105]=1;ram[122][106]=0;ram[122][107]=0;ram[122][108]=1;ram[122][109]=1;ram[122][110]=1;ram[122][111]=1;ram[122][112]=0;ram[122][113]=1;ram[122][114]=1;ram[122][115]=1;ram[122][116]=1;ram[122][117]=0;ram[122][118]=1;ram[122][119]=1;ram[122][120]=1;ram[122][121]=0;ram[122][122]=0;ram[122][123]=1;ram[122][124]=1;ram[122][125]=1;ram[122][126]=0;ram[122][127]=0;ram[122][128]=0;ram[122][129]=1;ram[122][130]=0;ram[122][131]=1;ram[122][132]=1;ram[122][133]=0;ram[122][134]=1;ram[122][135]=1;ram[122][136]=1;
        ram[123][0]=1;ram[123][1]=1;ram[123][2]=1;ram[123][3]=1;ram[123][4]=0;ram[123][5]=1;ram[123][6]=0;ram[123][7]=0;ram[123][8]=0;ram[123][9]=1;ram[123][10]=0;ram[123][11]=1;ram[123][12]=1;ram[123][13]=1;ram[123][14]=0;ram[123][15]=0;ram[123][16]=1;ram[123][17]=1;ram[123][18]=1;ram[123][19]=1;ram[123][20]=1;ram[123][21]=0;ram[123][22]=1;ram[123][23]=1;ram[123][24]=1;ram[123][25]=0;ram[123][26]=1;ram[123][27]=0;ram[123][28]=1;ram[123][29]=1;ram[123][30]=1;ram[123][31]=0;ram[123][32]=1;ram[123][33]=0;ram[123][34]=1;ram[123][35]=0;ram[123][36]=1;ram[123][37]=1;ram[123][38]=0;ram[123][39]=1;ram[123][40]=1;ram[123][41]=0;ram[123][42]=1;ram[123][43]=1;ram[123][44]=1;ram[123][45]=0;ram[123][46]=1;ram[123][47]=1;ram[123][48]=1;ram[123][49]=0;ram[123][50]=0;ram[123][51]=1;ram[123][52]=1;ram[123][53]=1;ram[123][54]=1;ram[123][55]=0;ram[123][56]=0;ram[123][57]=1;ram[123][58]=1;ram[123][59]=0;ram[123][60]=1;ram[123][61]=1;ram[123][62]=1;ram[123][63]=1;ram[123][64]=1;ram[123][65]=1;ram[123][66]=1;ram[123][67]=0;ram[123][68]=1;ram[123][69]=0;ram[123][70]=1;ram[123][71]=1;ram[123][72]=0;ram[123][73]=0;ram[123][74]=0;ram[123][75]=0;ram[123][76]=0;ram[123][77]=0;ram[123][78]=1;ram[123][79]=0;ram[123][80]=1;ram[123][81]=1;ram[123][82]=0;ram[123][83]=1;ram[123][84]=1;ram[123][85]=1;ram[123][86]=0;ram[123][87]=1;ram[123][88]=0;ram[123][89]=1;ram[123][90]=1;ram[123][91]=0;ram[123][92]=0;ram[123][93]=1;ram[123][94]=1;ram[123][95]=1;ram[123][96]=1;ram[123][97]=1;ram[123][98]=1;ram[123][99]=1;ram[123][100]=1;ram[123][101]=1;ram[123][102]=0;ram[123][103]=0;ram[123][104]=0;ram[123][105]=1;ram[123][106]=1;ram[123][107]=1;ram[123][108]=0;ram[123][109]=1;ram[123][110]=1;ram[123][111]=0;ram[123][112]=0;ram[123][113]=1;ram[123][114]=1;ram[123][115]=0;ram[123][116]=0;ram[123][117]=1;ram[123][118]=1;ram[123][119]=1;ram[123][120]=1;ram[123][121]=0;ram[123][122]=1;ram[123][123]=1;ram[123][124]=1;ram[123][125]=1;ram[123][126]=0;ram[123][127]=1;ram[123][128]=1;ram[123][129]=1;ram[123][130]=1;ram[123][131]=0;ram[123][132]=0;ram[123][133]=1;ram[123][134]=1;ram[123][135]=1;ram[123][136]=1;
        ram[124][0]=1;ram[124][1]=0;ram[124][2]=0;ram[124][3]=1;ram[124][4]=1;ram[124][5]=1;ram[124][6]=1;ram[124][7]=1;ram[124][8]=1;ram[124][9]=1;ram[124][10]=1;ram[124][11]=1;ram[124][12]=0;ram[124][13]=0;ram[124][14]=1;ram[124][15]=0;ram[124][16]=0;ram[124][17]=0;ram[124][18]=1;ram[124][19]=1;ram[124][20]=1;ram[124][21]=1;ram[124][22]=0;ram[124][23]=1;ram[124][24]=1;ram[124][25]=0;ram[124][26]=0;ram[124][27]=0;ram[124][28]=0;ram[124][29]=1;ram[124][30]=1;ram[124][31]=1;ram[124][32]=1;ram[124][33]=1;ram[124][34]=1;ram[124][35]=0;ram[124][36]=0;ram[124][37]=1;ram[124][38]=1;ram[124][39]=1;ram[124][40]=1;ram[124][41]=1;ram[124][42]=1;ram[124][43]=1;ram[124][44]=0;ram[124][45]=1;ram[124][46]=1;ram[124][47]=0;ram[124][48]=1;ram[124][49]=1;ram[124][50]=1;ram[124][51]=0;ram[124][52]=0;ram[124][53]=1;ram[124][54]=0;ram[124][55]=0;ram[124][56]=1;ram[124][57]=0;ram[124][58]=0;ram[124][59]=0;ram[124][60]=1;ram[124][61]=1;ram[124][62]=1;ram[124][63]=1;ram[124][64]=0;ram[124][65]=1;ram[124][66]=0;ram[124][67]=1;ram[124][68]=1;ram[124][69]=1;ram[124][70]=1;ram[124][71]=0;ram[124][72]=1;ram[124][73]=0;ram[124][74]=0;ram[124][75]=1;ram[124][76]=0;ram[124][77]=1;ram[124][78]=1;ram[124][79]=0;ram[124][80]=1;ram[124][81]=1;ram[124][82]=0;ram[124][83]=1;ram[124][84]=1;ram[124][85]=1;ram[124][86]=1;ram[124][87]=1;ram[124][88]=1;ram[124][89]=1;ram[124][90]=1;ram[124][91]=1;ram[124][92]=1;ram[124][93]=1;ram[124][94]=0;ram[124][95]=1;ram[124][96]=0;ram[124][97]=0;ram[124][98]=1;ram[124][99]=0;ram[124][100]=0;ram[124][101]=1;ram[124][102]=1;ram[124][103]=0;ram[124][104]=0;ram[124][105]=0;ram[124][106]=1;ram[124][107]=0;ram[124][108]=1;ram[124][109]=0;ram[124][110]=1;ram[124][111]=0;ram[124][112]=1;ram[124][113]=1;ram[124][114]=0;ram[124][115]=0;ram[124][116]=1;ram[124][117]=1;ram[124][118]=1;ram[124][119]=1;ram[124][120]=1;ram[124][121]=1;ram[124][122]=0;ram[124][123]=1;ram[124][124]=0;ram[124][125]=1;ram[124][126]=0;ram[124][127]=1;ram[124][128]=1;ram[124][129]=0;ram[124][130]=0;ram[124][131]=0;ram[124][132]=1;ram[124][133]=1;ram[124][134]=1;ram[124][135]=1;ram[124][136]=1;
        ram[125][0]=0;ram[125][1]=1;ram[125][2]=1;ram[125][3]=1;ram[125][4]=1;ram[125][5]=0;ram[125][6]=0;ram[125][7]=1;ram[125][8]=1;ram[125][9]=1;ram[125][10]=1;ram[125][11]=1;ram[125][12]=1;ram[125][13]=1;ram[125][14]=1;ram[125][15]=0;ram[125][16]=1;ram[125][17]=0;ram[125][18]=0;ram[125][19]=1;ram[125][20]=1;ram[125][21]=0;ram[125][22]=1;ram[125][23]=1;ram[125][24]=1;ram[125][25]=1;ram[125][26]=0;ram[125][27]=1;ram[125][28]=1;ram[125][29]=1;ram[125][30]=1;ram[125][31]=1;ram[125][32]=0;ram[125][33]=0;ram[125][34]=0;ram[125][35]=0;ram[125][36]=1;ram[125][37]=0;ram[125][38]=1;ram[125][39]=0;ram[125][40]=1;ram[125][41]=0;ram[125][42]=1;ram[125][43]=0;ram[125][44]=1;ram[125][45]=1;ram[125][46]=0;ram[125][47]=1;ram[125][48]=0;ram[125][49]=1;ram[125][50]=0;ram[125][51]=0;ram[125][52]=0;ram[125][53]=1;ram[125][54]=1;ram[125][55]=0;ram[125][56]=0;ram[125][57]=1;ram[125][58]=1;ram[125][59]=0;ram[125][60]=1;ram[125][61]=1;ram[125][62]=1;ram[125][63]=0;ram[125][64]=1;ram[125][65]=1;ram[125][66]=0;ram[125][67]=1;ram[125][68]=1;ram[125][69]=0;ram[125][70]=0;ram[125][71]=1;ram[125][72]=0;ram[125][73]=1;ram[125][74]=1;ram[125][75]=1;ram[125][76]=1;ram[125][77]=1;ram[125][78]=0;ram[125][79]=0;ram[125][80]=1;ram[125][81]=0;ram[125][82]=0;ram[125][83]=1;ram[125][84]=1;ram[125][85]=1;ram[125][86]=0;ram[125][87]=0;ram[125][88]=1;ram[125][89]=1;ram[125][90]=1;ram[125][91]=0;ram[125][92]=1;ram[125][93]=0;ram[125][94]=1;ram[125][95]=0;ram[125][96]=1;ram[125][97]=0;ram[125][98]=1;ram[125][99]=1;ram[125][100]=1;ram[125][101]=1;ram[125][102]=1;ram[125][103]=0;ram[125][104]=0;ram[125][105]=1;ram[125][106]=0;ram[125][107]=1;ram[125][108]=0;ram[125][109]=0;ram[125][110]=1;ram[125][111]=1;ram[125][112]=0;ram[125][113]=0;ram[125][114]=1;ram[125][115]=1;ram[125][116]=1;ram[125][117]=1;ram[125][118]=0;ram[125][119]=1;ram[125][120]=0;ram[125][121]=1;ram[125][122]=1;ram[125][123]=1;ram[125][124]=0;ram[125][125]=1;ram[125][126]=1;ram[125][127]=0;ram[125][128]=1;ram[125][129]=1;ram[125][130]=0;ram[125][131]=0;ram[125][132]=0;ram[125][133]=0;ram[125][134]=1;ram[125][135]=1;ram[125][136]=0;
        ram[126][0]=1;ram[126][1]=1;ram[126][2]=0;ram[126][3]=1;ram[126][4]=1;ram[126][5]=1;ram[126][6]=1;ram[126][7]=1;ram[126][8]=1;ram[126][9]=0;ram[126][10]=0;ram[126][11]=1;ram[126][12]=0;ram[126][13]=0;ram[126][14]=0;ram[126][15]=1;ram[126][16]=1;ram[126][17]=1;ram[126][18]=1;ram[126][19]=0;ram[126][20]=1;ram[126][21]=1;ram[126][22]=1;ram[126][23]=0;ram[126][24]=0;ram[126][25]=1;ram[126][26]=0;ram[126][27]=1;ram[126][28]=1;ram[126][29]=0;ram[126][30]=0;ram[126][31]=0;ram[126][32]=0;ram[126][33]=1;ram[126][34]=1;ram[126][35]=0;ram[126][36]=0;ram[126][37]=1;ram[126][38]=1;ram[126][39]=1;ram[126][40]=1;ram[126][41]=1;ram[126][42]=1;ram[126][43]=0;ram[126][44]=0;ram[126][45]=0;ram[126][46]=0;ram[126][47]=0;ram[126][48]=1;ram[126][49]=1;ram[126][50]=0;ram[126][51]=1;ram[126][52]=1;ram[126][53]=1;ram[126][54]=1;ram[126][55]=1;ram[126][56]=1;ram[126][57]=1;ram[126][58]=0;ram[126][59]=0;ram[126][60]=1;ram[126][61]=1;ram[126][62]=1;ram[126][63]=0;ram[126][64]=0;ram[126][65]=1;ram[126][66]=1;ram[126][67]=0;ram[126][68]=1;ram[126][69]=1;ram[126][70]=1;ram[126][71]=1;ram[126][72]=1;ram[126][73]=1;ram[126][74]=1;ram[126][75]=1;ram[126][76]=0;ram[126][77]=0;ram[126][78]=1;ram[126][79]=1;ram[126][80]=1;ram[126][81]=1;ram[126][82]=0;ram[126][83]=1;ram[126][84]=0;ram[126][85]=0;ram[126][86]=0;ram[126][87]=1;ram[126][88]=0;ram[126][89]=1;ram[126][90]=1;ram[126][91]=1;ram[126][92]=1;ram[126][93]=1;ram[126][94]=0;ram[126][95]=1;ram[126][96]=0;ram[126][97]=1;ram[126][98]=1;ram[126][99]=1;ram[126][100]=1;ram[126][101]=0;ram[126][102]=1;ram[126][103]=0;ram[126][104]=1;ram[126][105]=1;ram[126][106]=1;ram[126][107]=1;ram[126][108]=0;ram[126][109]=1;ram[126][110]=0;ram[126][111]=0;ram[126][112]=1;ram[126][113]=0;ram[126][114]=0;ram[126][115]=1;ram[126][116]=1;ram[126][117]=1;ram[126][118]=1;ram[126][119]=1;ram[126][120]=0;ram[126][121]=1;ram[126][122]=1;ram[126][123]=1;ram[126][124]=0;ram[126][125]=0;ram[126][126]=0;ram[126][127]=0;ram[126][128]=1;ram[126][129]=0;ram[126][130]=1;ram[126][131]=1;ram[126][132]=1;ram[126][133]=0;ram[126][134]=1;ram[126][135]=1;ram[126][136]=0;
        ram[127][0]=0;ram[127][1]=1;ram[127][2]=0;ram[127][3]=1;ram[127][4]=0;ram[127][5]=1;ram[127][6]=1;ram[127][7]=1;ram[127][8]=0;ram[127][9]=1;ram[127][10]=1;ram[127][11]=1;ram[127][12]=1;ram[127][13]=1;ram[127][14]=1;ram[127][15]=1;ram[127][16]=1;ram[127][17]=1;ram[127][18]=1;ram[127][19]=0;ram[127][20]=0;ram[127][21]=1;ram[127][22]=0;ram[127][23]=1;ram[127][24]=1;ram[127][25]=0;ram[127][26]=1;ram[127][27]=1;ram[127][28]=0;ram[127][29]=1;ram[127][30]=0;ram[127][31]=0;ram[127][32]=0;ram[127][33]=1;ram[127][34]=1;ram[127][35]=0;ram[127][36]=1;ram[127][37]=1;ram[127][38]=0;ram[127][39]=1;ram[127][40]=1;ram[127][41]=0;ram[127][42]=1;ram[127][43]=1;ram[127][44]=1;ram[127][45]=1;ram[127][46]=1;ram[127][47]=0;ram[127][48]=0;ram[127][49]=1;ram[127][50]=1;ram[127][51]=1;ram[127][52]=0;ram[127][53]=1;ram[127][54]=1;ram[127][55]=1;ram[127][56]=1;ram[127][57]=1;ram[127][58]=1;ram[127][59]=1;ram[127][60]=1;ram[127][61]=1;ram[127][62]=0;ram[127][63]=1;ram[127][64]=0;ram[127][65]=0;ram[127][66]=1;ram[127][67]=1;ram[127][68]=0;ram[127][69]=1;ram[127][70]=0;ram[127][71]=0;ram[127][72]=1;ram[127][73]=1;ram[127][74]=1;ram[127][75]=1;ram[127][76]=1;ram[127][77]=1;ram[127][78]=0;ram[127][79]=0;ram[127][80]=1;ram[127][81]=1;ram[127][82]=0;ram[127][83]=1;ram[127][84]=0;ram[127][85]=0;ram[127][86]=0;ram[127][87]=0;ram[127][88]=1;ram[127][89]=1;ram[127][90]=1;ram[127][91]=1;ram[127][92]=0;ram[127][93]=1;ram[127][94]=0;ram[127][95]=0;ram[127][96]=1;ram[127][97]=1;ram[127][98]=1;ram[127][99]=1;ram[127][100]=1;ram[127][101]=0;ram[127][102]=0;ram[127][103]=1;ram[127][104]=1;ram[127][105]=1;ram[127][106]=0;ram[127][107]=1;ram[127][108]=1;ram[127][109]=1;ram[127][110]=1;ram[127][111]=1;ram[127][112]=1;ram[127][113]=0;ram[127][114]=1;ram[127][115]=0;ram[127][116]=0;ram[127][117]=1;ram[127][118]=1;ram[127][119]=1;ram[127][120]=0;ram[127][121]=1;ram[127][122]=1;ram[127][123]=0;ram[127][124]=0;ram[127][125]=1;ram[127][126]=0;ram[127][127]=1;ram[127][128]=0;ram[127][129]=0;ram[127][130]=1;ram[127][131]=1;ram[127][132]=1;ram[127][133]=0;ram[127][134]=0;ram[127][135]=1;ram[127][136]=1;
        ram[128][0]=0;ram[128][1]=1;ram[128][2]=1;ram[128][3]=1;ram[128][4]=1;ram[128][5]=0;ram[128][6]=1;ram[128][7]=0;ram[128][8]=1;ram[128][9]=1;ram[128][10]=0;ram[128][11]=0;ram[128][12]=1;ram[128][13]=1;ram[128][14]=1;ram[128][15]=0;ram[128][16]=1;ram[128][17]=1;ram[128][18]=1;ram[128][19]=1;ram[128][20]=1;ram[128][21]=1;ram[128][22]=1;ram[128][23]=1;ram[128][24]=1;ram[128][25]=0;ram[128][26]=1;ram[128][27]=0;ram[128][28]=1;ram[128][29]=1;ram[128][30]=1;ram[128][31]=1;ram[128][32]=0;ram[128][33]=1;ram[128][34]=0;ram[128][35]=1;ram[128][36]=0;ram[128][37]=1;ram[128][38]=1;ram[128][39]=0;ram[128][40]=1;ram[128][41]=0;ram[128][42]=0;ram[128][43]=0;ram[128][44]=0;ram[128][45]=0;ram[128][46]=0;ram[128][47]=0;ram[128][48]=0;ram[128][49]=1;ram[128][50]=0;ram[128][51]=1;ram[128][52]=1;ram[128][53]=0;ram[128][54]=0;ram[128][55]=0;ram[128][56]=1;ram[128][57]=1;ram[128][58]=1;ram[128][59]=1;ram[128][60]=0;ram[128][61]=1;ram[128][62]=0;ram[128][63]=0;ram[128][64]=0;ram[128][65]=1;ram[128][66]=1;ram[128][67]=1;ram[128][68]=1;ram[128][69]=0;ram[128][70]=0;ram[128][71]=1;ram[128][72]=0;ram[128][73]=1;ram[128][74]=0;ram[128][75]=0;ram[128][76]=1;ram[128][77]=0;ram[128][78]=1;ram[128][79]=1;ram[128][80]=1;ram[128][81]=1;ram[128][82]=1;ram[128][83]=1;ram[128][84]=1;ram[128][85]=1;ram[128][86]=0;ram[128][87]=1;ram[128][88]=1;ram[128][89]=1;ram[128][90]=1;ram[128][91]=0;ram[128][92]=1;ram[128][93]=1;ram[128][94]=1;ram[128][95]=1;ram[128][96]=0;ram[128][97]=1;ram[128][98]=0;ram[128][99]=1;ram[128][100]=1;ram[128][101]=1;ram[128][102]=1;ram[128][103]=0;ram[128][104]=1;ram[128][105]=0;ram[128][106]=1;ram[128][107]=0;ram[128][108]=1;ram[128][109]=1;ram[128][110]=0;ram[128][111]=0;ram[128][112]=0;ram[128][113]=1;ram[128][114]=1;ram[128][115]=0;ram[128][116]=1;ram[128][117]=1;ram[128][118]=0;ram[128][119]=0;ram[128][120]=0;ram[128][121]=0;ram[128][122]=1;ram[128][123]=1;ram[128][124]=1;ram[128][125]=1;ram[128][126]=0;ram[128][127]=1;ram[128][128]=1;ram[128][129]=0;ram[128][130]=0;ram[128][131]=0;ram[128][132]=1;ram[128][133]=0;ram[128][134]=0;ram[128][135]=1;ram[128][136]=0;
        ram[129][0]=1;ram[129][1]=0;ram[129][2]=0;ram[129][3]=1;ram[129][4]=1;ram[129][5]=1;ram[129][6]=0;ram[129][7]=0;ram[129][8]=1;ram[129][9]=1;ram[129][10]=0;ram[129][11]=0;ram[129][12]=1;ram[129][13]=1;ram[129][14]=1;ram[129][15]=1;ram[129][16]=0;ram[129][17]=1;ram[129][18]=1;ram[129][19]=1;ram[129][20]=0;ram[129][21]=0;ram[129][22]=0;ram[129][23]=1;ram[129][24]=1;ram[129][25]=0;ram[129][26]=1;ram[129][27]=1;ram[129][28]=0;ram[129][29]=1;ram[129][30]=1;ram[129][31]=1;ram[129][32]=0;ram[129][33]=1;ram[129][34]=0;ram[129][35]=0;ram[129][36]=1;ram[129][37]=1;ram[129][38]=1;ram[129][39]=1;ram[129][40]=1;ram[129][41]=1;ram[129][42]=0;ram[129][43]=0;ram[129][44]=0;ram[129][45]=1;ram[129][46]=1;ram[129][47]=1;ram[129][48]=1;ram[129][49]=1;ram[129][50]=0;ram[129][51]=1;ram[129][52]=0;ram[129][53]=0;ram[129][54]=1;ram[129][55]=1;ram[129][56]=1;ram[129][57]=1;ram[129][58]=0;ram[129][59]=1;ram[129][60]=1;ram[129][61]=1;ram[129][62]=1;ram[129][63]=0;ram[129][64]=1;ram[129][65]=1;ram[129][66]=1;ram[129][67]=0;ram[129][68]=1;ram[129][69]=1;ram[129][70]=1;ram[129][71]=1;ram[129][72]=1;ram[129][73]=0;ram[129][74]=0;ram[129][75]=1;ram[129][76]=1;ram[129][77]=1;ram[129][78]=1;ram[129][79]=0;ram[129][80]=1;ram[129][81]=1;ram[129][82]=1;ram[129][83]=1;ram[129][84]=1;ram[129][85]=0;ram[129][86]=1;ram[129][87]=1;ram[129][88]=1;ram[129][89]=0;ram[129][90]=0;ram[129][91]=1;ram[129][92]=1;ram[129][93]=0;ram[129][94]=0;ram[129][95]=0;ram[129][96]=0;ram[129][97]=1;ram[129][98]=1;ram[129][99]=1;ram[129][100]=1;ram[129][101]=0;ram[129][102]=1;ram[129][103]=1;ram[129][104]=0;ram[129][105]=1;ram[129][106]=1;ram[129][107]=1;ram[129][108]=1;ram[129][109]=1;ram[129][110]=1;ram[129][111]=1;ram[129][112]=0;ram[129][113]=0;ram[129][114]=1;ram[129][115]=1;ram[129][116]=0;ram[129][117]=1;ram[129][118]=1;ram[129][119]=1;ram[129][120]=0;ram[129][121]=1;ram[129][122]=1;ram[129][123]=0;ram[129][124]=0;ram[129][125]=0;ram[129][126]=0;ram[129][127]=1;ram[129][128]=0;ram[129][129]=0;ram[129][130]=0;ram[129][131]=1;ram[129][132]=1;ram[129][133]=1;ram[129][134]=1;ram[129][135]=1;ram[129][136]=0;
        ram[130][0]=0;ram[130][1]=1;ram[130][2]=0;ram[130][3]=0;ram[130][4]=1;ram[130][5]=1;ram[130][6]=0;ram[130][7]=1;ram[130][8]=0;ram[130][9]=0;ram[130][10]=1;ram[130][11]=0;ram[130][12]=1;ram[130][13]=1;ram[130][14]=1;ram[130][15]=0;ram[130][16]=1;ram[130][17]=0;ram[130][18]=0;ram[130][19]=0;ram[130][20]=1;ram[130][21]=1;ram[130][22]=1;ram[130][23]=1;ram[130][24]=1;ram[130][25]=1;ram[130][26]=0;ram[130][27]=1;ram[130][28]=1;ram[130][29]=1;ram[130][30]=0;ram[130][31]=1;ram[130][32]=1;ram[130][33]=1;ram[130][34]=1;ram[130][35]=0;ram[130][36]=1;ram[130][37]=0;ram[130][38]=1;ram[130][39]=0;ram[130][40]=0;ram[130][41]=1;ram[130][42]=1;ram[130][43]=1;ram[130][44]=1;ram[130][45]=1;ram[130][46]=1;ram[130][47]=1;ram[130][48]=1;ram[130][49]=0;ram[130][50]=0;ram[130][51]=1;ram[130][52]=0;ram[130][53]=1;ram[130][54]=1;ram[130][55]=0;ram[130][56]=1;ram[130][57]=1;ram[130][58]=0;ram[130][59]=1;ram[130][60]=0;ram[130][61]=1;ram[130][62]=1;ram[130][63]=0;ram[130][64]=0;ram[130][65]=0;ram[130][66]=0;ram[130][67]=1;ram[130][68]=1;ram[130][69]=1;ram[130][70]=1;ram[130][71]=1;ram[130][72]=1;ram[130][73]=1;ram[130][74]=0;ram[130][75]=1;ram[130][76]=1;ram[130][77]=1;ram[130][78]=0;ram[130][79]=0;ram[130][80]=1;ram[130][81]=0;ram[130][82]=1;ram[130][83]=0;ram[130][84]=1;ram[130][85]=1;ram[130][86]=1;ram[130][87]=1;ram[130][88]=1;ram[130][89]=1;ram[130][90]=1;ram[130][91]=1;ram[130][92]=0;ram[130][93]=0;ram[130][94]=1;ram[130][95]=1;ram[130][96]=1;ram[130][97]=0;ram[130][98]=1;ram[130][99]=1;ram[130][100]=1;ram[130][101]=1;ram[130][102]=0;ram[130][103]=0;ram[130][104]=1;ram[130][105]=1;ram[130][106]=1;ram[130][107]=1;ram[130][108]=1;ram[130][109]=1;ram[130][110]=0;ram[130][111]=1;ram[130][112]=1;ram[130][113]=1;ram[130][114]=1;ram[130][115]=0;ram[130][116]=0;ram[130][117]=1;ram[130][118]=0;ram[130][119]=0;ram[130][120]=1;ram[130][121]=1;ram[130][122]=1;ram[130][123]=0;ram[130][124]=1;ram[130][125]=0;ram[130][126]=0;ram[130][127]=1;ram[130][128]=1;ram[130][129]=1;ram[130][130]=0;ram[130][131]=0;ram[130][132]=0;ram[130][133]=1;ram[130][134]=0;ram[130][135]=0;ram[130][136]=1;
        ram[131][0]=1;ram[131][1]=1;ram[131][2]=0;ram[131][3]=1;ram[131][4]=0;ram[131][5]=0;ram[131][6]=1;ram[131][7]=1;ram[131][8]=1;ram[131][9]=1;ram[131][10]=0;ram[131][11]=1;ram[131][12]=1;ram[131][13]=1;ram[131][14]=0;ram[131][15]=0;ram[131][16]=1;ram[131][17]=1;ram[131][18]=1;ram[131][19]=0;ram[131][20]=1;ram[131][21]=1;ram[131][22]=1;ram[131][23]=0;ram[131][24]=0;ram[131][25]=1;ram[131][26]=0;ram[131][27]=1;ram[131][28]=1;ram[131][29]=1;ram[131][30]=1;ram[131][31]=1;ram[131][32]=0;ram[131][33]=0;ram[131][34]=0;ram[131][35]=1;ram[131][36]=1;ram[131][37]=1;ram[131][38]=1;ram[131][39]=1;ram[131][40]=1;ram[131][41]=1;ram[131][42]=0;ram[131][43]=0;ram[131][44]=0;ram[131][45]=1;ram[131][46]=1;ram[131][47]=1;ram[131][48]=1;ram[131][49]=1;ram[131][50]=1;ram[131][51]=1;ram[131][52]=0;ram[131][53]=0;ram[131][54]=0;ram[131][55]=0;ram[131][56]=0;ram[131][57]=1;ram[131][58]=1;ram[131][59]=0;ram[131][60]=1;ram[131][61]=1;ram[131][62]=1;ram[131][63]=0;ram[131][64]=1;ram[131][65]=1;ram[131][66]=1;ram[131][67]=0;ram[131][68]=1;ram[131][69]=0;ram[131][70]=1;ram[131][71]=1;ram[131][72]=0;ram[131][73]=1;ram[131][74]=1;ram[131][75]=0;ram[131][76]=1;ram[131][77]=0;ram[131][78]=1;ram[131][79]=1;ram[131][80]=1;ram[131][81]=1;ram[131][82]=1;ram[131][83]=1;ram[131][84]=1;ram[131][85]=0;ram[131][86]=1;ram[131][87]=1;ram[131][88]=1;ram[131][89]=1;ram[131][90]=1;ram[131][91]=1;ram[131][92]=0;ram[131][93]=1;ram[131][94]=1;ram[131][95]=0;ram[131][96]=1;ram[131][97]=1;ram[131][98]=0;ram[131][99]=1;ram[131][100]=0;ram[131][101]=1;ram[131][102]=1;ram[131][103]=0;ram[131][104]=0;ram[131][105]=1;ram[131][106]=0;ram[131][107]=1;ram[131][108]=1;ram[131][109]=1;ram[131][110]=1;ram[131][111]=0;ram[131][112]=1;ram[131][113]=0;ram[131][114]=1;ram[131][115]=0;ram[131][116]=1;ram[131][117]=1;ram[131][118]=1;ram[131][119]=1;ram[131][120]=1;ram[131][121]=1;ram[131][122]=1;ram[131][123]=0;ram[131][124]=1;ram[131][125]=1;ram[131][126]=1;ram[131][127]=1;ram[131][128]=1;ram[131][129]=0;ram[131][130]=0;ram[131][131]=1;ram[131][132]=0;ram[131][133]=0;ram[131][134]=0;ram[131][135]=1;ram[131][136]=1;
        ram[132][0]=1;ram[132][1]=1;ram[132][2]=0;ram[132][3]=0;ram[132][4]=0;ram[132][5]=1;ram[132][6]=0;ram[132][7]=0;ram[132][8]=1;ram[132][9]=0;ram[132][10]=0;ram[132][11]=0;ram[132][12]=0;ram[132][13]=1;ram[132][14]=0;ram[132][15]=1;ram[132][16]=1;ram[132][17]=0;ram[132][18]=1;ram[132][19]=1;ram[132][20]=0;ram[132][21]=1;ram[132][22]=1;ram[132][23]=1;ram[132][24]=1;ram[132][25]=1;ram[132][26]=1;ram[132][27]=1;ram[132][28]=1;ram[132][29]=0;ram[132][30]=0;ram[132][31]=0;ram[132][32]=1;ram[132][33]=1;ram[132][34]=1;ram[132][35]=1;ram[132][36]=1;ram[132][37]=0;ram[132][38]=1;ram[132][39]=1;ram[132][40]=1;ram[132][41]=0;ram[132][42]=1;ram[132][43]=0;ram[132][44]=1;ram[132][45]=1;ram[132][46]=1;ram[132][47]=1;ram[132][48]=0;ram[132][49]=1;ram[132][50]=0;ram[132][51]=0;ram[132][52]=1;ram[132][53]=0;ram[132][54]=0;ram[132][55]=1;ram[132][56]=1;ram[132][57]=1;ram[132][58]=1;ram[132][59]=1;ram[132][60]=0;ram[132][61]=1;ram[132][62]=0;ram[132][63]=0;ram[132][64]=0;ram[132][65]=1;ram[132][66]=1;ram[132][67]=1;ram[132][68]=0;ram[132][69]=0;ram[132][70]=0;ram[132][71]=0;ram[132][72]=1;ram[132][73]=1;ram[132][74]=1;ram[132][75]=1;ram[132][76]=1;ram[132][77]=1;ram[132][78]=1;ram[132][79]=1;ram[132][80]=1;ram[132][81]=0;ram[132][82]=0;ram[132][83]=1;ram[132][84]=1;ram[132][85]=1;ram[132][86]=0;ram[132][87]=1;ram[132][88]=0;ram[132][89]=0;ram[132][90]=1;ram[132][91]=1;ram[132][92]=1;ram[132][93]=1;ram[132][94]=1;ram[132][95]=1;ram[132][96]=1;ram[132][97]=1;ram[132][98]=1;ram[132][99]=1;ram[132][100]=1;ram[132][101]=1;ram[132][102]=1;ram[132][103]=1;ram[132][104]=0;ram[132][105]=0;ram[132][106]=1;ram[132][107]=1;ram[132][108]=1;ram[132][109]=0;ram[132][110]=1;ram[132][111]=1;ram[132][112]=1;ram[132][113]=0;ram[132][114]=1;ram[132][115]=1;ram[132][116]=1;ram[132][117]=1;ram[132][118]=1;ram[132][119]=0;ram[132][120]=1;ram[132][121]=1;ram[132][122]=0;ram[132][123]=0;ram[132][124]=0;ram[132][125]=0;ram[132][126]=1;ram[132][127]=0;ram[132][128]=1;ram[132][129]=0;ram[132][130]=1;ram[132][131]=1;ram[132][132]=1;ram[132][133]=1;ram[132][134]=1;ram[132][135]=1;ram[132][136]=1;
        ram[133][0]=0;ram[133][1]=1;ram[133][2]=0;ram[133][3]=1;ram[133][4]=1;ram[133][5]=1;ram[133][6]=0;ram[133][7]=0;ram[133][8]=1;ram[133][9]=1;ram[133][10]=1;ram[133][11]=0;ram[133][12]=0;ram[133][13]=1;ram[133][14]=1;ram[133][15]=1;ram[133][16]=1;ram[133][17]=0;ram[133][18]=0;ram[133][19]=1;ram[133][20]=1;ram[133][21]=1;ram[133][22]=1;ram[133][23]=1;ram[133][24]=1;ram[133][25]=0;ram[133][26]=1;ram[133][27]=1;ram[133][28]=0;ram[133][29]=1;ram[133][30]=1;ram[133][31]=1;ram[133][32]=1;ram[133][33]=0;ram[133][34]=1;ram[133][35]=0;ram[133][36]=1;ram[133][37]=1;ram[133][38]=1;ram[133][39]=1;ram[133][40]=1;ram[133][41]=1;ram[133][42]=0;ram[133][43]=1;ram[133][44]=1;ram[133][45]=1;ram[133][46]=0;ram[133][47]=1;ram[133][48]=1;ram[133][49]=1;ram[133][50]=1;ram[133][51]=1;ram[133][52]=0;ram[133][53]=1;ram[133][54]=0;ram[133][55]=1;ram[133][56]=1;ram[133][57]=0;ram[133][58]=1;ram[133][59]=1;ram[133][60]=0;ram[133][61]=1;ram[133][62]=1;ram[133][63]=1;ram[133][64]=1;ram[133][65]=0;ram[133][66]=1;ram[133][67]=1;ram[133][68]=1;ram[133][69]=1;ram[133][70]=0;ram[133][71]=1;ram[133][72]=0;ram[133][73]=1;ram[133][74]=1;ram[133][75]=1;ram[133][76]=1;ram[133][77]=1;ram[133][78]=1;ram[133][79]=1;ram[133][80]=1;ram[133][81]=1;ram[133][82]=0;ram[133][83]=0;ram[133][84]=0;ram[133][85]=0;ram[133][86]=1;ram[133][87]=0;ram[133][88]=0;ram[133][89]=1;ram[133][90]=1;ram[133][91]=0;ram[133][92]=0;ram[133][93]=1;ram[133][94]=1;ram[133][95]=1;ram[133][96]=1;ram[133][97]=0;ram[133][98]=0;ram[133][99]=0;ram[133][100]=1;ram[133][101]=1;ram[133][102]=0;ram[133][103]=0;ram[133][104]=1;ram[133][105]=0;ram[133][106]=1;ram[133][107]=1;ram[133][108]=1;ram[133][109]=1;ram[133][110]=1;ram[133][111]=0;ram[133][112]=1;ram[133][113]=1;ram[133][114]=1;ram[133][115]=0;ram[133][116]=0;ram[133][117]=1;ram[133][118]=1;ram[133][119]=1;ram[133][120]=1;ram[133][121]=1;ram[133][122]=1;ram[133][123]=1;ram[133][124]=1;ram[133][125]=1;ram[133][126]=1;ram[133][127]=1;ram[133][128]=0;ram[133][129]=0;ram[133][130]=1;ram[133][131]=1;ram[133][132]=1;ram[133][133]=0;ram[133][134]=0;ram[133][135]=1;ram[133][136]=0;
        ram[134][0]=1;ram[134][1]=1;ram[134][2]=1;ram[134][3]=1;ram[134][4]=0;ram[134][5]=1;ram[134][6]=0;ram[134][7]=0;ram[134][8]=0;ram[134][9]=1;ram[134][10]=1;ram[134][11]=0;ram[134][12]=1;ram[134][13]=0;ram[134][14]=1;ram[134][15]=0;ram[134][16]=1;ram[134][17]=0;ram[134][18]=0;ram[134][19]=1;ram[134][20]=1;ram[134][21]=0;ram[134][22]=1;ram[134][23]=1;ram[134][24]=1;ram[134][25]=1;ram[134][26]=1;ram[134][27]=1;ram[134][28]=0;ram[134][29]=1;ram[134][30]=0;ram[134][31]=0;ram[134][32]=1;ram[134][33]=1;ram[134][34]=1;ram[134][35]=1;ram[134][36]=1;ram[134][37]=0;ram[134][38]=1;ram[134][39]=0;ram[134][40]=0;ram[134][41]=0;ram[134][42]=0;ram[134][43]=1;ram[134][44]=1;ram[134][45]=1;ram[134][46]=1;ram[134][47]=1;ram[134][48]=1;ram[134][49]=1;ram[134][50]=1;ram[134][51]=0;ram[134][52]=1;ram[134][53]=1;ram[134][54]=1;ram[134][55]=1;ram[134][56]=0;ram[134][57]=1;ram[134][58]=0;ram[134][59]=1;ram[134][60]=1;ram[134][61]=0;ram[134][62]=1;ram[134][63]=1;ram[134][64]=1;ram[134][65]=1;ram[134][66]=0;ram[134][67]=1;ram[134][68]=1;ram[134][69]=0;ram[134][70]=1;ram[134][71]=0;ram[134][72]=1;ram[134][73]=1;ram[134][74]=1;ram[134][75]=1;ram[134][76]=1;ram[134][77]=1;ram[134][78]=0;ram[134][79]=1;ram[134][80]=1;ram[134][81]=1;ram[134][82]=1;ram[134][83]=1;ram[134][84]=1;ram[134][85]=1;ram[134][86]=0;ram[134][87]=0;ram[134][88]=1;ram[134][89]=0;ram[134][90]=1;ram[134][91]=1;ram[134][92]=1;ram[134][93]=1;ram[134][94]=0;ram[134][95]=1;ram[134][96]=1;ram[134][97]=0;ram[134][98]=0;ram[134][99]=1;ram[134][100]=1;ram[134][101]=0;ram[134][102]=1;ram[134][103]=1;ram[134][104]=0;ram[134][105]=0;ram[134][106]=1;ram[134][107]=1;ram[134][108]=0;ram[134][109]=0;ram[134][110]=0;ram[134][111]=1;ram[134][112]=1;ram[134][113]=1;ram[134][114]=0;ram[134][115]=1;ram[134][116]=1;ram[134][117]=1;ram[134][118]=0;ram[134][119]=1;ram[134][120]=0;ram[134][121]=1;ram[134][122]=0;ram[134][123]=0;ram[134][124]=1;ram[134][125]=0;ram[134][126]=1;ram[134][127]=1;ram[134][128]=1;ram[134][129]=0;ram[134][130]=1;ram[134][131]=1;ram[134][132]=1;ram[134][133]=1;ram[134][134]=1;ram[134][135]=0;ram[134][136]=1;
        ram[135][0]=0;ram[135][1]=1;ram[135][2]=1;ram[135][3]=0;ram[135][4]=1;ram[135][5]=1;ram[135][6]=0;ram[135][7]=1;ram[135][8]=1;ram[135][9]=1;ram[135][10]=1;ram[135][11]=1;ram[135][12]=0;ram[135][13]=0;ram[135][14]=1;ram[135][15]=1;ram[135][16]=0;ram[135][17]=1;ram[135][18]=1;ram[135][19]=1;ram[135][20]=1;ram[135][21]=0;ram[135][22]=1;ram[135][23]=0;ram[135][24]=1;ram[135][25]=1;ram[135][26]=1;ram[135][27]=1;ram[135][28]=0;ram[135][29]=1;ram[135][30]=1;ram[135][31]=1;ram[135][32]=1;ram[135][33]=0;ram[135][34]=1;ram[135][35]=1;ram[135][36]=0;ram[135][37]=1;ram[135][38]=1;ram[135][39]=0;ram[135][40]=1;ram[135][41]=1;ram[135][42]=1;ram[135][43]=1;ram[135][44]=1;ram[135][45]=0;ram[135][46]=0;ram[135][47]=0;ram[135][48]=1;ram[135][49]=1;ram[135][50]=1;ram[135][51]=0;ram[135][52]=0;ram[135][53]=0;ram[135][54]=1;ram[135][55]=1;ram[135][56]=0;ram[135][57]=1;ram[135][58]=0;ram[135][59]=0;ram[135][60]=1;ram[135][61]=1;ram[135][62]=1;ram[135][63]=0;ram[135][64]=1;ram[135][65]=1;ram[135][66]=1;ram[135][67]=1;ram[135][68]=1;ram[135][69]=1;ram[135][70]=1;ram[135][71]=1;ram[135][72]=1;ram[135][73]=1;ram[135][74]=0;ram[135][75]=1;ram[135][76]=1;ram[135][77]=0;ram[135][78]=0;ram[135][79]=1;ram[135][80]=1;ram[135][81]=0;ram[135][82]=1;ram[135][83]=1;ram[135][84]=1;ram[135][85]=1;ram[135][86]=1;ram[135][87]=0;ram[135][88]=0;ram[135][89]=0;ram[135][90]=1;ram[135][91]=0;ram[135][92]=0;ram[135][93]=0;ram[135][94]=1;ram[135][95]=1;ram[135][96]=1;ram[135][97]=1;ram[135][98]=1;ram[135][99]=1;ram[135][100]=1;ram[135][101]=0;ram[135][102]=0;ram[135][103]=0;ram[135][104]=0;ram[135][105]=1;ram[135][106]=1;ram[135][107]=1;ram[135][108]=0;ram[135][109]=1;ram[135][110]=1;ram[135][111]=0;ram[135][112]=0;ram[135][113]=1;ram[135][114]=1;ram[135][115]=1;ram[135][116]=1;ram[135][117]=0;ram[135][118]=0;ram[135][119]=1;ram[135][120]=0;ram[135][121]=0;ram[135][122]=1;ram[135][123]=0;ram[135][124]=0;ram[135][125]=1;ram[135][126]=1;ram[135][127]=1;ram[135][128]=0;ram[135][129]=1;ram[135][130]=1;ram[135][131]=0;ram[135][132]=1;ram[135][133]=1;ram[135][134]=1;ram[135][135]=0;ram[135][136]=0;
        ram[136][0]=1;ram[136][1]=1;ram[136][2]=0;ram[136][3]=0;ram[136][4]=0;ram[136][5]=0;ram[136][6]=0;ram[136][7]=0;ram[136][8]=0;ram[136][9]=0;ram[136][10]=1;ram[136][11]=0;ram[136][12]=1;ram[136][13]=1;ram[136][14]=1;ram[136][15]=1;ram[136][16]=0;ram[136][17]=1;ram[136][18]=1;ram[136][19]=0;ram[136][20]=0;ram[136][21]=0;ram[136][22]=1;ram[136][23]=1;ram[136][24]=0;ram[136][25]=0;ram[136][26]=0;ram[136][27]=0;ram[136][28]=1;ram[136][29]=1;ram[136][30]=1;ram[136][31]=0;ram[136][32]=0;ram[136][33]=0;ram[136][34]=1;ram[136][35]=0;ram[136][36]=1;ram[136][37]=0;ram[136][38]=1;ram[136][39]=0;ram[136][40]=0;ram[136][41]=1;ram[136][42]=1;ram[136][43]=1;ram[136][44]=0;ram[136][45]=0;ram[136][46]=1;ram[136][47]=1;ram[136][48]=0;ram[136][49]=1;ram[136][50]=1;ram[136][51]=1;ram[136][52]=0;ram[136][53]=1;ram[136][54]=1;ram[136][55]=0;ram[136][56]=0;ram[136][57]=1;ram[136][58]=0;ram[136][59]=0;ram[136][60]=1;ram[136][61]=1;ram[136][62]=1;ram[136][63]=1;ram[136][64]=1;ram[136][65]=0;ram[136][66]=1;ram[136][67]=1;ram[136][68]=0;ram[136][69]=1;ram[136][70]=1;ram[136][71]=0;ram[136][72]=0;ram[136][73]=0;ram[136][74]=0;ram[136][75]=1;ram[136][76]=0;ram[136][77]=1;ram[136][78]=0;ram[136][79]=0;ram[136][80]=0;ram[136][81]=0;ram[136][82]=1;ram[136][83]=1;ram[136][84]=1;ram[136][85]=0;ram[136][86]=1;ram[136][87]=1;ram[136][88]=1;ram[136][89]=1;ram[136][90]=0;ram[136][91]=0;ram[136][92]=1;ram[136][93]=1;ram[136][94]=1;ram[136][95]=0;ram[136][96]=1;ram[136][97]=1;ram[136][98]=1;ram[136][99]=1;ram[136][100]=1;ram[136][101]=0;ram[136][102]=0;ram[136][103]=0;ram[136][104]=1;ram[136][105]=1;ram[136][106]=1;ram[136][107]=1;ram[136][108]=1;ram[136][109]=1;ram[136][110]=1;ram[136][111]=0;ram[136][112]=1;ram[136][113]=1;ram[136][114]=1;ram[136][115]=1;ram[136][116]=1;ram[136][117]=1;ram[136][118]=1;ram[136][119]=1;ram[136][120]=1;ram[136][121]=1;ram[136][122]=1;ram[136][123]=0;ram[136][124]=0;ram[136][125]=0;ram[136][126]=1;ram[136][127]=1;ram[136][128]=1;ram[136][129]=1;ram[136][130]=0;ram[136][131]=1;ram[136][132]=0;ram[136][133]=0;ram[136][134]=1;ram[136][135]=1;ram[136][136]=0;

        sum<=0;
    end
    
    genvar i;
    genvar j;
    generate
        for(i=0;i<size;i=i+1)
        begin: row
            for(j=0;j<size;j=j+1)
            begin: column
            
                if( (i==0 && (j==0 || j==size-1)) || (i==size-1 && (j==0 || j==size-1)) )
                begin: i_j_zero
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else sumram[i][j]=1;
                    end
                end
                
                else if(i==0)
                begin: i_zero
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else if (ram[i][j-1]+ram[i][j+1]+ram[i+1][j-1]+ram[i+1][j]+ram[i+1][j+1]<4)sumram[i][j]=1;
                        else sumram[i][j]=0;
                    end
                end
                
                else if(i==size-1)
                begin: i_end
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else if (ram[i][j-1]+ram[i][j+1]+ram[i-1][j-1]+ram[i-1][j]+ram[i-1][j+1]<4)sumram[i][j]=1;
                        else sumram[i][j]=0;
                    end
                end
                
                else if(j==0)
                begin: j_zero
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else if (ram[i-1][j]+ram[i-1][j+1]+ram[i][j+1]+ram[i+1][j]+ram[i+1][j+1]<4)sumram[i][j]=1;
                        else sumram[i][j]=0;
                    end
                end
                
                else if(j==size-1)
                begin: j_end
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else if (ram[i-1][j-1]+ram[i-1][j]+ram[i][j-1]+ram[i+1][j-1]+ram[i+1][j]<4)sumram[i][j]=1;
                        else sumram[i][j]=0;
                    end
                end
                
                else
                begin: normal
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else if (ram[i-1][j-1]+ram[i-1][j]+ram[i-1][j+1]+ram[i][j-1]+ram[i][j+1]+ram[i+1][j-1]+ram[i+1][j]+ram[i+1][j+1]<4)sumram[i][j]=1;
                        else sumram[i][j]=0;
                    end
                end
            end
        end
    endgenerate
    
    wire [8:0]sumcache[size-1:0];
    assign sumcache[0]=sumram[0][0]+sumram[0][1]+sumram[0][2]+sumram[0][3]+sumram[0][4]+sumram[0][5]+sumram[0][6]+sumram[0][7]+sumram[0][8]+sumram[0][9]+sumram[0][10]+sumram[0][11]+sumram[0][12]+sumram[0][13]+sumram[0][14]+sumram[0][15]+sumram[0][16]+sumram[0][17]+sumram[0][18]+sumram[0][19]+sumram[0][20]+sumram[0][21]+sumram[0][22]+sumram[0][23]+sumram[0][24]+sumram[0][25]+sumram[0][26]+sumram[0][27]+sumram[0][28]+sumram[0][29]+sumram[0][30]+sumram[0][31]+sumram[0][32]+sumram[0][33]+sumram[0][34]+sumram[0][35]+sumram[0][36]+sumram[0][37]+sumram[0][38]+sumram[0][39]+sumram[0][40]+sumram[0][41]+sumram[0][42]+sumram[0][43]+sumram[0][44]+sumram[0][45]+sumram[0][46]+sumram[0][47]+sumram[0][48]+sumram[0][49]+sumram[0][50]+sumram[0][51]+sumram[0][52]+sumram[0][53]+sumram[0][54]+sumram[0][55]+sumram[0][56]+sumram[0][57]+sumram[0][58]+sumram[0][59]+sumram[0][60]+sumram[0][61]+sumram[0][62]+sumram[0][63]+sumram[0][64]+sumram[0][65]+sumram[0][66]+sumram[0][67]+sumram[0][68]+sumram[0][69]+sumram[0][70]+sumram[0][71]+sumram[0][72]+sumram[0][73]+sumram[0][74]+sumram[0][75]+sumram[0][76]+sumram[0][77]+sumram[0][78]+sumram[0][79]+sumram[0][80]+sumram[0][81]+sumram[0][82]+sumram[0][83]+sumram[0][84]+sumram[0][85]+sumram[0][86]+sumram[0][87]+sumram[0][88]+sumram[0][89]+sumram[0][90]+sumram[0][91]+sumram[0][92]+sumram[0][93]+sumram[0][94]+sumram[0][95]+sumram[0][96]+sumram[0][97]+sumram[0][98]+sumram[0][99]+sumram[0][100]+sumram[0][101]+sumram[0][102]+sumram[0][103]+sumram[0][104]+sumram[0][105]+sumram[0][106]+sumram[0][107]+sumram[0][108]+sumram[0][109]+sumram[0][110]+sumram[0][111]+sumram[0][112]+sumram[0][113]+sumram[0][114]+sumram[0][115]+sumram[0][116]+sumram[0][117]+sumram[0][118]+sumram[0][119]+sumram[0][120]+sumram[0][121]+sumram[0][122]+sumram[0][123]+sumram[0][124]+sumram[0][125]+sumram[0][126]+sumram[0][127]+sumram[0][128]+sumram[0][129]+sumram[0][130]+sumram[0][131]+sumram[0][132]+sumram[0][133]+sumram[0][134]+sumram[0][135]+sumram[0][136];
    assign sumcache[1]=sumram[1][0]+sumram[1][1]+sumram[1][2]+sumram[1][3]+sumram[1][4]+sumram[1][5]+sumram[1][6]+sumram[1][7]+sumram[1][8]+sumram[1][9]+sumram[1][10]+sumram[1][11]+sumram[1][12]+sumram[1][13]+sumram[1][14]+sumram[1][15]+sumram[1][16]+sumram[1][17]+sumram[1][18]+sumram[1][19]+sumram[1][20]+sumram[1][21]+sumram[1][22]+sumram[1][23]+sumram[1][24]+sumram[1][25]+sumram[1][26]+sumram[1][27]+sumram[1][28]+sumram[1][29]+sumram[1][30]+sumram[1][31]+sumram[1][32]+sumram[1][33]+sumram[1][34]+sumram[1][35]+sumram[1][36]+sumram[1][37]+sumram[1][38]+sumram[1][39]+sumram[1][40]+sumram[1][41]+sumram[1][42]+sumram[1][43]+sumram[1][44]+sumram[1][45]+sumram[1][46]+sumram[1][47]+sumram[1][48]+sumram[1][49]+sumram[1][50]+sumram[1][51]+sumram[1][52]+sumram[1][53]+sumram[1][54]+sumram[1][55]+sumram[1][56]+sumram[1][57]+sumram[1][58]+sumram[1][59]+sumram[1][60]+sumram[1][61]+sumram[1][62]+sumram[1][63]+sumram[1][64]+sumram[1][65]+sumram[1][66]+sumram[1][67]+sumram[1][68]+sumram[1][69]+sumram[1][70]+sumram[1][71]+sumram[1][72]+sumram[1][73]+sumram[1][74]+sumram[1][75]+sumram[1][76]+sumram[1][77]+sumram[1][78]+sumram[1][79]+sumram[1][80]+sumram[1][81]+sumram[1][82]+sumram[1][83]+sumram[1][84]+sumram[1][85]+sumram[1][86]+sumram[1][87]+sumram[1][88]+sumram[1][89]+sumram[1][90]+sumram[1][91]+sumram[1][92]+sumram[1][93]+sumram[1][94]+sumram[1][95]+sumram[1][96]+sumram[1][97]+sumram[1][98]+sumram[1][99]+sumram[1][100]+sumram[1][101]+sumram[1][102]+sumram[1][103]+sumram[1][104]+sumram[1][105]+sumram[1][106]+sumram[1][107]+sumram[1][108]+sumram[1][109]+sumram[1][110]+sumram[1][111]+sumram[1][112]+sumram[1][113]+sumram[1][114]+sumram[1][115]+sumram[1][116]+sumram[1][117]+sumram[1][118]+sumram[1][119]+sumram[1][120]+sumram[1][121]+sumram[1][122]+sumram[1][123]+sumram[1][124]+sumram[1][125]+sumram[1][126]+sumram[1][127]+sumram[1][128]+sumram[1][129]+sumram[1][130]+sumram[1][131]+sumram[1][132]+sumram[1][133]+sumram[1][134]+sumram[1][135]+sumram[1][136];
    assign sumcache[2]=sumram[2][0]+sumram[2][1]+sumram[2][2]+sumram[2][3]+sumram[2][4]+sumram[2][5]+sumram[2][6]+sumram[2][7]+sumram[2][8]+sumram[2][9]+sumram[2][10]+sumram[2][11]+sumram[2][12]+sumram[2][13]+sumram[2][14]+sumram[2][15]+sumram[2][16]+sumram[2][17]+sumram[2][18]+sumram[2][19]+sumram[2][20]+sumram[2][21]+sumram[2][22]+sumram[2][23]+sumram[2][24]+sumram[2][25]+sumram[2][26]+sumram[2][27]+sumram[2][28]+sumram[2][29]+sumram[2][30]+sumram[2][31]+sumram[2][32]+sumram[2][33]+sumram[2][34]+sumram[2][35]+sumram[2][36]+sumram[2][37]+sumram[2][38]+sumram[2][39]+sumram[2][40]+sumram[2][41]+sumram[2][42]+sumram[2][43]+sumram[2][44]+sumram[2][45]+sumram[2][46]+sumram[2][47]+sumram[2][48]+sumram[2][49]+sumram[2][50]+sumram[2][51]+sumram[2][52]+sumram[2][53]+sumram[2][54]+sumram[2][55]+sumram[2][56]+sumram[2][57]+sumram[2][58]+sumram[2][59]+sumram[2][60]+sumram[2][61]+sumram[2][62]+sumram[2][63]+sumram[2][64]+sumram[2][65]+sumram[2][66]+sumram[2][67]+sumram[2][68]+sumram[2][69]+sumram[2][70]+sumram[2][71]+sumram[2][72]+sumram[2][73]+sumram[2][74]+sumram[2][75]+sumram[2][76]+sumram[2][77]+sumram[2][78]+sumram[2][79]+sumram[2][80]+sumram[2][81]+sumram[2][82]+sumram[2][83]+sumram[2][84]+sumram[2][85]+sumram[2][86]+sumram[2][87]+sumram[2][88]+sumram[2][89]+sumram[2][90]+sumram[2][91]+sumram[2][92]+sumram[2][93]+sumram[2][94]+sumram[2][95]+sumram[2][96]+sumram[2][97]+sumram[2][98]+sumram[2][99]+sumram[2][100]+sumram[2][101]+sumram[2][102]+sumram[2][103]+sumram[2][104]+sumram[2][105]+sumram[2][106]+sumram[2][107]+sumram[2][108]+sumram[2][109]+sumram[2][110]+sumram[2][111]+sumram[2][112]+sumram[2][113]+sumram[2][114]+sumram[2][115]+sumram[2][116]+sumram[2][117]+sumram[2][118]+sumram[2][119]+sumram[2][120]+sumram[2][121]+sumram[2][122]+sumram[2][123]+sumram[2][124]+sumram[2][125]+sumram[2][126]+sumram[2][127]+sumram[2][128]+sumram[2][129]+sumram[2][130]+sumram[2][131]+sumram[2][132]+sumram[2][133]+sumram[2][134]+sumram[2][135]+sumram[2][136];
    assign sumcache[3]=sumram[3][0]+sumram[3][1]+sumram[3][2]+sumram[3][3]+sumram[3][4]+sumram[3][5]+sumram[3][6]+sumram[3][7]+sumram[3][8]+sumram[3][9]+sumram[3][10]+sumram[3][11]+sumram[3][12]+sumram[3][13]+sumram[3][14]+sumram[3][15]+sumram[3][16]+sumram[3][17]+sumram[3][18]+sumram[3][19]+sumram[3][20]+sumram[3][21]+sumram[3][22]+sumram[3][23]+sumram[3][24]+sumram[3][25]+sumram[3][26]+sumram[3][27]+sumram[3][28]+sumram[3][29]+sumram[3][30]+sumram[3][31]+sumram[3][32]+sumram[3][33]+sumram[3][34]+sumram[3][35]+sumram[3][36]+sumram[3][37]+sumram[3][38]+sumram[3][39]+sumram[3][40]+sumram[3][41]+sumram[3][42]+sumram[3][43]+sumram[3][44]+sumram[3][45]+sumram[3][46]+sumram[3][47]+sumram[3][48]+sumram[3][49]+sumram[3][50]+sumram[3][51]+sumram[3][52]+sumram[3][53]+sumram[3][54]+sumram[3][55]+sumram[3][56]+sumram[3][57]+sumram[3][58]+sumram[3][59]+sumram[3][60]+sumram[3][61]+sumram[3][62]+sumram[3][63]+sumram[3][64]+sumram[3][65]+sumram[3][66]+sumram[3][67]+sumram[3][68]+sumram[3][69]+sumram[3][70]+sumram[3][71]+sumram[3][72]+sumram[3][73]+sumram[3][74]+sumram[3][75]+sumram[3][76]+sumram[3][77]+sumram[3][78]+sumram[3][79]+sumram[3][80]+sumram[3][81]+sumram[3][82]+sumram[3][83]+sumram[3][84]+sumram[3][85]+sumram[3][86]+sumram[3][87]+sumram[3][88]+sumram[3][89]+sumram[3][90]+sumram[3][91]+sumram[3][92]+sumram[3][93]+sumram[3][94]+sumram[3][95]+sumram[3][96]+sumram[3][97]+sumram[3][98]+sumram[3][99]+sumram[3][100]+sumram[3][101]+sumram[3][102]+sumram[3][103]+sumram[3][104]+sumram[3][105]+sumram[3][106]+sumram[3][107]+sumram[3][108]+sumram[3][109]+sumram[3][110]+sumram[3][111]+sumram[3][112]+sumram[3][113]+sumram[3][114]+sumram[3][115]+sumram[3][116]+sumram[3][117]+sumram[3][118]+sumram[3][119]+sumram[3][120]+sumram[3][121]+sumram[3][122]+sumram[3][123]+sumram[3][124]+sumram[3][125]+sumram[3][126]+sumram[3][127]+sumram[3][128]+sumram[3][129]+sumram[3][130]+sumram[3][131]+sumram[3][132]+sumram[3][133]+sumram[3][134]+sumram[3][135]+sumram[3][136];
    assign sumcache[4]=sumram[4][0]+sumram[4][1]+sumram[4][2]+sumram[4][3]+sumram[4][4]+sumram[4][5]+sumram[4][6]+sumram[4][7]+sumram[4][8]+sumram[4][9]+sumram[4][10]+sumram[4][11]+sumram[4][12]+sumram[4][13]+sumram[4][14]+sumram[4][15]+sumram[4][16]+sumram[4][17]+sumram[4][18]+sumram[4][19]+sumram[4][20]+sumram[4][21]+sumram[4][22]+sumram[4][23]+sumram[4][24]+sumram[4][25]+sumram[4][26]+sumram[4][27]+sumram[4][28]+sumram[4][29]+sumram[4][30]+sumram[4][31]+sumram[4][32]+sumram[4][33]+sumram[4][34]+sumram[4][35]+sumram[4][36]+sumram[4][37]+sumram[4][38]+sumram[4][39]+sumram[4][40]+sumram[4][41]+sumram[4][42]+sumram[4][43]+sumram[4][44]+sumram[4][45]+sumram[4][46]+sumram[4][47]+sumram[4][48]+sumram[4][49]+sumram[4][50]+sumram[4][51]+sumram[4][52]+sumram[4][53]+sumram[4][54]+sumram[4][55]+sumram[4][56]+sumram[4][57]+sumram[4][58]+sumram[4][59]+sumram[4][60]+sumram[4][61]+sumram[4][62]+sumram[4][63]+sumram[4][64]+sumram[4][65]+sumram[4][66]+sumram[4][67]+sumram[4][68]+sumram[4][69]+sumram[4][70]+sumram[4][71]+sumram[4][72]+sumram[4][73]+sumram[4][74]+sumram[4][75]+sumram[4][76]+sumram[4][77]+sumram[4][78]+sumram[4][79]+sumram[4][80]+sumram[4][81]+sumram[4][82]+sumram[4][83]+sumram[4][84]+sumram[4][85]+sumram[4][86]+sumram[4][87]+sumram[4][88]+sumram[4][89]+sumram[4][90]+sumram[4][91]+sumram[4][92]+sumram[4][93]+sumram[4][94]+sumram[4][95]+sumram[4][96]+sumram[4][97]+sumram[4][98]+sumram[4][99]+sumram[4][100]+sumram[4][101]+sumram[4][102]+sumram[4][103]+sumram[4][104]+sumram[4][105]+sumram[4][106]+sumram[4][107]+sumram[4][108]+sumram[4][109]+sumram[4][110]+sumram[4][111]+sumram[4][112]+sumram[4][113]+sumram[4][114]+sumram[4][115]+sumram[4][116]+sumram[4][117]+sumram[4][118]+sumram[4][119]+sumram[4][120]+sumram[4][121]+sumram[4][122]+sumram[4][123]+sumram[4][124]+sumram[4][125]+sumram[4][126]+sumram[4][127]+sumram[4][128]+sumram[4][129]+sumram[4][130]+sumram[4][131]+sumram[4][132]+sumram[4][133]+sumram[4][134]+sumram[4][135]+sumram[4][136];
    assign sumcache[5]=sumram[5][0]+sumram[5][1]+sumram[5][2]+sumram[5][3]+sumram[5][4]+sumram[5][5]+sumram[5][6]+sumram[5][7]+sumram[5][8]+sumram[5][9]+sumram[5][10]+sumram[5][11]+sumram[5][12]+sumram[5][13]+sumram[5][14]+sumram[5][15]+sumram[5][16]+sumram[5][17]+sumram[5][18]+sumram[5][19]+sumram[5][20]+sumram[5][21]+sumram[5][22]+sumram[5][23]+sumram[5][24]+sumram[5][25]+sumram[5][26]+sumram[5][27]+sumram[5][28]+sumram[5][29]+sumram[5][30]+sumram[5][31]+sumram[5][32]+sumram[5][33]+sumram[5][34]+sumram[5][35]+sumram[5][36]+sumram[5][37]+sumram[5][38]+sumram[5][39]+sumram[5][40]+sumram[5][41]+sumram[5][42]+sumram[5][43]+sumram[5][44]+sumram[5][45]+sumram[5][46]+sumram[5][47]+sumram[5][48]+sumram[5][49]+sumram[5][50]+sumram[5][51]+sumram[5][52]+sumram[5][53]+sumram[5][54]+sumram[5][55]+sumram[5][56]+sumram[5][57]+sumram[5][58]+sumram[5][59]+sumram[5][60]+sumram[5][61]+sumram[5][62]+sumram[5][63]+sumram[5][64]+sumram[5][65]+sumram[5][66]+sumram[5][67]+sumram[5][68]+sumram[5][69]+sumram[5][70]+sumram[5][71]+sumram[5][72]+sumram[5][73]+sumram[5][74]+sumram[5][75]+sumram[5][76]+sumram[5][77]+sumram[5][78]+sumram[5][79]+sumram[5][80]+sumram[5][81]+sumram[5][82]+sumram[5][83]+sumram[5][84]+sumram[5][85]+sumram[5][86]+sumram[5][87]+sumram[5][88]+sumram[5][89]+sumram[5][90]+sumram[5][91]+sumram[5][92]+sumram[5][93]+sumram[5][94]+sumram[5][95]+sumram[5][96]+sumram[5][97]+sumram[5][98]+sumram[5][99]+sumram[5][100]+sumram[5][101]+sumram[5][102]+sumram[5][103]+sumram[5][104]+sumram[5][105]+sumram[5][106]+sumram[5][107]+sumram[5][108]+sumram[5][109]+sumram[5][110]+sumram[5][111]+sumram[5][112]+sumram[5][113]+sumram[5][114]+sumram[5][115]+sumram[5][116]+sumram[5][117]+sumram[5][118]+sumram[5][119]+sumram[5][120]+sumram[5][121]+sumram[5][122]+sumram[5][123]+sumram[5][124]+sumram[5][125]+sumram[5][126]+sumram[5][127]+sumram[5][128]+sumram[5][129]+sumram[5][130]+sumram[5][131]+sumram[5][132]+sumram[5][133]+sumram[5][134]+sumram[5][135]+sumram[5][136];
    assign sumcache[6]=sumram[6][0]+sumram[6][1]+sumram[6][2]+sumram[6][3]+sumram[6][4]+sumram[6][5]+sumram[6][6]+sumram[6][7]+sumram[6][8]+sumram[6][9]+sumram[6][10]+sumram[6][11]+sumram[6][12]+sumram[6][13]+sumram[6][14]+sumram[6][15]+sumram[6][16]+sumram[6][17]+sumram[6][18]+sumram[6][19]+sumram[6][20]+sumram[6][21]+sumram[6][22]+sumram[6][23]+sumram[6][24]+sumram[6][25]+sumram[6][26]+sumram[6][27]+sumram[6][28]+sumram[6][29]+sumram[6][30]+sumram[6][31]+sumram[6][32]+sumram[6][33]+sumram[6][34]+sumram[6][35]+sumram[6][36]+sumram[6][37]+sumram[6][38]+sumram[6][39]+sumram[6][40]+sumram[6][41]+sumram[6][42]+sumram[6][43]+sumram[6][44]+sumram[6][45]+sumram[6][46]+sumram[6][47]+sumram[6][48]+sumram[6][49]+sumram[6][50]+sumram[6][51]+sumram[6][52]+sumram[6][53]+sumram[6][54]+sumram[6][55]+sumram[6][56]+sumram[6][57]+sumram[6][58]+sumram[6][59]+sumram[6][60]+sumram[6][61]+sumram[6][62]+sumram[6][63]+sumram[6][64]+sumram[6][65]+sumram[6][66]+sumram[6][67]+sumram[6][68]+sumram[6][69]+sumram[6][70]+sumram[6][71]+sumram[6][72]+sumram[6][73]+sumram[6][74]+sumram[6][75]+sumram[6][76]+sumram[6][77]+sumram[6][78]+sumram[6][79]+sumram[6][80]+sumram[6][81]+sumram[6][82]+sumram[6][83]+sumram[6][84]+sumram[6][85]+sumram[6][86]+sumram[6][87]+sumram[6][88]+sumram[6][89]+sumram[6][90]+sumram[6][91]+sumram[6][92]+sumram[6][93]+sumram[6][94]+sumram[6][95]+sumram[6][96]+sumram[6][97]+sumram[6][98]+sumram[6][99]+sumram[6][100]+sumram[6][101]+sumram[6][102]+sumram[6][103]+sumram[6][104]+sumram[6][105]+sumram[6][106]+sumram[6][107]+sumram[6][108]+sumram[6][109]+sumram[6][110]+sumram[6][111]+sumram[6][112]+sumram[6][113]+sumram[6][114]+sumram[6][115]+sumram[6][116]+sumram[6][117]+sumram[6][118]+sumram[6][119]+sumram[6][120]+sumram[6][121]+sumram[6][122]+sumram[6][123]+sumram[6][124]+sumram[6][125]+sumram[6][126]+sumram[6][127]+sumram[6][128]+sumram[6][129]+sumram[6][130]+sumram[6][131]+sumram[6][132]+sumram[6][133]+sumram[6][134]+sumram[6][135]+sumram[6][136];
    assign sumcache[7]=sumram[7][0]+sumram[7][1]+sumram[7][2]+sumram[7][3]+sumram[7][4]+sumram[7][5]+sumram[7][6]+sumram[7][7]+sumram[7][8]+sumram[7][9]+sumram[7][10]+sumram[7][11]+sumram[7][12]+sumram[7][13]+sumram[7][14]+sumram[7][15]+sumram[7][16]+sumram[7][17]+sumram[7][18]+sumram[7][19]+sumram[7][20]+sumram[7][21]+sumram[7][22]+sumram[7][23]+sumram[7][24]+sumram[7][25]+sumram[7][26]+sumram[7][27]+sumram[7][28]+sumram[7][29]+sumram[7][30]+sumram[7][31]+sumram[7][32]+sumram[7][33]+sumram[7][34]+sumram[7][35]+sumram[7][36]+sumram[7][37]+sumram[7][38]+sumram[7][39]+sumram[7][40]+sumram[7][41]+sumram[7][42]+sumram[7][43]+sumram[7][44]+sumram[7][45]+sumram[7][46]+sumram[7][47]+sumram[7][48]+sumram[7][49]+sumram[7][50]+sumram[7][51]+sumram[7][52]+sumram[7][53]+sumram[7][54]+sumram[7][55]+sumram[7][56]+sumram[7][57]+sumram[7][58]+sumram[7][59]+sumram[7][60]+sumram[7][61]+sumram[7][62]+sumram[7][63]+sumram[7][64]+sumram[7][65]+sumram[7][66]+sumram[7][67]+sumram[7][68]+sumram[7][69]+sumram[7][70]+sumram[7][71]+sumram[7][72]+sumram[7][73]+sumram[7][74]+sumram[7][75]+sumram[7][76]+sumram[7][77]+sumram[7][78]+sumram[7][79]+sumram[7][80]+sumram[7][81]+sumram[7][82]+sumram[7][83]+sumram[7][84]+sumram[7][85]+sumram[7][86]+sumram[7][87]+sumram[7][88]+sumram[7][89]+sumram[7][90]+sumram[7][91]+sumram[7][92]+sumram[7][93]+sumram[7][94]+sumram[7][95]+sumram[7][96]+sumram[7][97]+sumram[7][98]+sumram[7][99]+sumram[7][100]+sumram[7][101]+sumram[7][102]+sumram[7][103]+sumram[7][104]+sumram[7][105]+sumram[7][106]+sumram[7][107]+sumram[7][108]+sumram[7][109]+sumram[7][110]+sumram[7][111]+sumram[7][112]+sumram[7][113]+sumram[7][114]+sumram[7][115]+sumram[7][116]+sumram[7][117]+sumram[7][118]+sumram[7][119]+sumram[7][120]+sumram[7][121]+sumram[7][122]+sumram[7][123]+sumram[7][124]+sumram[7][125]+sumram[7][126]+sumram[7][127]+sumram[7][128]+sumram[7][129]+sumram[7][130]+sumram[7][131]+sumram[7][132]+sumram[7][133]+sumram[7][134]+sumram[7][135]+sumram[7][136];
    assign sumcache[8]=sumram[8][0]+sumram[8][1]+sumram[8][2]+sumram[8][3]+sumram[8][4]+sumram[8][5]+sumram[8][6]+sumram[8][7]+sumram[8][8]+sumram[8][9]+sumram[8][10]+sumram[8][11]+sumram[8][12]+sumram[8][13]+sumram[8][14]+sumram[8][15]+sumram[8][16]+sumram[8][17]+sumram[8][18]+sumram[8][19]+sumram[8][20]+sumram[8][21]+sumram[8][22]+sumram[8][23]+sumram[8][24]+sumram[8][25]+sumram[8][26]+sumram[8][27]+sumram[8][28]+sumram[8][29]+sumram[8][30]+sumram[8][31]+sumram[8][32]+sumram[8][33]+sumram[8][34]+sumram[8][35]+sumram[8][36]+sumram[8][37]+sumram[8][38]+sumram[8][39]+sumram[8][40]+sumram[8][41]+sumram[8][42]+sumram[8][43]+sumram[8][44]+sumram[8][45]+sumram[8][46]+sumram[8][47]+sumram[8][48]+sumram[8][49]+sumram[8][50]+sumram[8][51]+sumram[8][52]+sumram[8][53]+sumram[8][54]+sumram[8][55]+sumram[8][56]+sumram[8][57]+sumram[8][58]+sumram[8][59]+sumram[8][60]+sumram[8][61]+sumram[8][62]+sumram[8][63]+sumram[8][64]+sumram[8][65]+sumram[8][66]+sumram[8][67]+sumram[8][68]+sumram[8][69]+sumram[8][70]+sumram[8][71]+sumram[8][72]+sumram[8][73]+sumram[8][74]+sumram[8][75]+sumram[8][76]+sumram[8][77]+sumram[8][78]+sumram[8][79]+sumram[8][80]+sumram[8][81]+sumram[8][82]+sumram[8][83]+sumram[8][84]+sumram[8][85]+sumram[8][86]+sumram[8][87]+sumram[8][88]+sumram[8][89]+sumram[8][90]+sumram[8][91]+sumram[8][92]+sumram[8][93]+sumram[8][94]+sumram[8][95]+sumram[8][96]+sumram[8][97]+sumram[8][98]+sumram[8][99]+sumram[8][100]+sumram[8][101]+sumram[8][102]+sumram[8][103]+sumram[8][104]+sumram[8][105]+sumram[8][106]+sumram[8][107]+sumram[8][108]+sumram[8][109]+sumram[8][110]+sumram[8][111]+sumram[8][112]+sumram[8][113]+sumram[8][114]+sumram[8][115]+sumram[8][116]+sumram[8][117]+sumram[8][118]+sumram[8][119]+sumram[8][120]+sumram[8][121]+sumram[8][122]+sumram[8][123]+sumram[8][124]+sumram[8][125]+sumram[8][126]+sumram[8][127]+sumram[8][128]+sumram[8][129]+sumram[8][130]+sumram[8][131]+sumram[8][132]+sumram[8][133]+sumram[8][134]+sumram[8][135]+sumram[8][136];
    assign sumcache[9]=sumram[9][0]+sumram[9][1]+sumram[9][2]+sumram[9][3]+sumram[9][4]+sumram[9][5]+sumram[9][6]+sumram[9][7]+sumram[9][8]+sumram[9][9]+sumram[9][10]+sumram[9][11]+sumram[9][12]+sumram[9][13]+sumram[9][14]+sumram[9][15]+sumram[9][16]+sumram[9][17]+sumram[9][18]+sumram[9][19]+sumram[9][20]+sumram[9][21]+sumram[9][22]+sumram[9][23]+sumram[9][24]+sumram[9][25]+sumram[9][26]+sumram[9][27]+sumram[9][28]+sumram[9][29]+sumram[9][30]+sumram[9][31]+sumram[9][32]+sumram[9][33]+sumram[9][34]+sumram[9][35]+sumram[9][36]+sumram[9][37]+sumram[9][38]+sumram[9][39]+sumram[9][40]+sumram[9][41]+sumram[9][42]+sumram[9][43]+sumram[9][44]+sumram[9][45]+sumram[9][46]+sumram[9][47]+sumram[9][48]+sumram[9][49]+sumram[9][50]+sumram[9][51]+sumram[9][52]+sumram[9][53]+sumram[9][54]+sumram[9][55]+sumram[9][56]+sumram[9][57]+sumram[9][58]+sumram[9][59]+sumram[9][60]+sumram[9][61]+sumram[9][62]+sumram[9][63]+sumram[9][64]+sumram[9][65]+sumram[9][66]+sumram[9][67]+sumram[9][68]+sumram[9][69]+sumram[9][70]+sumram[9][71]+sumram[9][72]+sumram[9][73]+sumram[9][74]+sumram[9][75]+sumram[9][76]+sumram[9][77]+sumram[9][78]+sumram[9][79]+sumram[9][80]+sumram[9][81]+sumram[9][82]+sumram[9][83]+sumram[9][84]+sumram[9][85]+sumram[9][86]+sumram[9][87]+sumram[9][88]+sumram[9][89]+sumram[9][90]+sumram[9][91]+sumram[9][92]+sumram[9][93]+sumram[9][94]+sumram[9][95]+sumram[9][96]+sumram[9][97]+sumram[9][98]+sumram[9][99]+sumram[9][100]+sumram[9][101]+sumram[9][102]+sumram[9][103]+sumram[9][104]+sumram[9][105]+sumram[9][106]+sumram[9][107]+sumram[9][108]+sumram[9][109]+sumram[9][110]+sumram[9][111]+sumram[9][112]+sumram[9][113]+sumram[9][114]+sumram[9][115]+sumram[9][116]+sumram[9][117]+sumram[9][118]+sumram[9][119]+sumram[9][120]+sumram[9][121]+sumram[9][122]+sumram[9][123]+sumram[9][124]+sumram[9][125]+sumram[9][126]+sumram[9][127]+sumram[9][128]+sumram[9][129]+sumram[9][130]+sumram[9][131]+sumram[9][132]+sumram[9][133]+sumram[9][134]+sumram[9][135]+sumram[9][136];
    assign sumcache[10]=sumram[10][0]+sumram[10][1]+sumram[10][2]+sumram[10][3]+sumram[10][4]+sumram[10][5]+sumram[10][6]+sumram[10][7]+sumram[10][8]+sumram[10][9]+sumram[10][10]+sumram[10][11]+sumram[10][12]+sumram[10][13]+sumram[10][14]+sumram[10][15]+sumram[10][16]+sumram[10][17]+sumram[10][18]+sumram[10][19]+sumram[10][20]+sumram[10][21]+sumram[10][22]+sumram[10][23]+sumram[10][24]+sumram[10][25]+sumram[10][26]+sumram[10][27]+sumram[10][28]+sumram[10][29]+sumram[10][30]+sumram[10][31]+sumram[10][32]+sumram[10][33]+sumram[10][34]+sumram[10][35]+sumram[10][36]+sumram[10][37]+sumram[10][38]+sumram[10][39]+sumram[10][40]+sumram[10][41]+sumram[10][42]+sumram[10][43]+sumram[10][44]+sumram[10][45]+sumram[10][46]+sumram[10][47]+sumram[10][48]+sumram[10][49]+sumram[10][50]+sumram[10][51]+sumram[10][52]+sumram[10][53]+sumram[10][54]+sumram[10][55]+sumram[10][56]+sumram[10][57]+sumram[10][58]+sumram[10][59]+sumram[10][60]+sumram[10][61]+sumram[10][62]+sumram[10][63]+sumram[10][64]+sumram[10][65]+sumram[10][66]+sumram[10][67]+sumram[10][68]+sumram[10][69]+sumram[10][70]+sumram[10][71]+sumram[10][72]+sumram[10][73]+sumram[10][74]+sumram[10][75]+sumram[10][76]+sumram[10][77]+sumram[10][78]+sumram[10][79]+sumram[10][80]+sumram[10][81]+sumram[10][82]+sumram[10][83]+sumram[10][84]+sumram[10][85]+sumram[10][86]+sumram[10][87]+sumram[10][88]+sumram[10][89]+sumram[10][90]+sumram[10][91]+sumram[10][92]+sumram[10][93]+sumram[10][94]+sumram[10][95]+sumram[10][96]+sumram[10][97]+sumram[10][98]+sumram[10][99]+sumram[10][100]+sumram[10][101]+sumram[10][102]+sumram[10][103]+sumram[10][104]+sumram[10][105]+sumram[10][106]+sumram[10][107]+sumram[10][108]+sumram[10][109]+sumram[10][110]+sumram[10][111]+sumram[10][112]+sumram[10][113]+sumram[10][114]+sumram[10][115]+sumram[10][116]+sumram[10][117]+sumram[10][118]+sumram[10][119]+sumram[10][120]+sumram[10][121]+sumram[10][122]+sumram[10][123]+sumram[10][124]+sumram[10][125]+sumram[10][126]+sumram[10][127]+sumram[10][128]+sumram[10][129]+sumram[10][130]+sumram[10][131]+sumram[10][132]+sumram[10][133]+sumram[10][134]+sumram[10][135]+sumram[10][136];
    assign sumcache[11]=sumram[11][0]+sumram[11][1]+sumram[11][2]+sumram[11][3]+sumram[11][4]+sumram[11][5]+sumram[11][6]+sumram[11][7]+sumram[11][8]+sumram[11][9]+sumram[11][10]+sumram[11][11]+sumram[11][12]+sumram[11][13]+sumram[11][14]+sumram[11][15]+sumram[11][16]+sumram[11][17]+sumram[11][18]+sumram[11][19]+sumram[11][20]+sumram[11][21]+sumram[11][22]+sumram[11][23]+sumram[11][24]+sumram[11][25]+sumram[11][26]+sumram[11][27]+sumram[11][28]+sumram[11][29]+sumram[11][30]+sumram[11][31]+sumram[11][32]+sumram[11][33]+sumram[11][34]+sumram[11][35]+sumram[11][36]+sumram[11][37]+sumram[11][38]+sumram[11][39]+sumram[11][40]+sumram[11][41]+sumram[11][42]+sumram[11][43]+sumram[11][44]+sumram[11][45]+sumram[11][46]+sumram[11][47]+sumram[11][48]+sumram[11][49]+sumram[11][50]+sumram[11][51]+sumram[11][52]+sumram[11][53]+sumram[11][54]+sumram[11][55]+sumram[11][56]+sumram[11][57]+sumram[11][58]+sumram[11][59]+sumram[11][60]+sumram[11][61]+sumram[11][62]+sumram[11][63]+sumram[11][64]+sumram[11][65]+sumram[11][66]+sumram[11][67]+sumram[11][68]+sumram[11][69]+sumram[11][70]+sumram[11][71]+sumram[11][72]+sumram[11][73]+sumram[11][74]+sumram[11][75]+sumram[11][76]+sumram[11][77]+sumram[11][78]+sumram[11][79]+sumram[11][80]+sumram[11][81]+sumram[11][82]+sumram[11][83]+sumram[11][84]+sumram[11][85]+sumram[11][86]+sumram[11][87]+sumram[11][88]+sumram[11][89]+sumram[11][90]+sumram[11][91]+sumram[11][92]+sumram[11][93]+sumram[11][94]+sumram[11][95]+sumram[11][96]+sumram[11][97]+sumram[11][98]+sumram[11][99]+sumram[11][100]+sumram[11][101]+sumram[11][102]+sumram[11][103]+sumram[11][104]+sumram[11][105]+sumram[11][106]+sumram[11][107]+sumram[11][108]+sumram[11][109]+sumram[11][110]+sumram[11][111]+sumram[11][112]+sumram[11][113]+sumram[11][114]+sumram[11][115]+sumram[11][116]+sumram[11][117]+sumram[11][118]+sumram[11][119]+sumram[11][120]+sumram[11][121]+sumram[11][122]+sumram[11][123]+sumram[11][124]+sumram[11][125]+sumram[11][126]+sumram[11][127]+sumram[11][128]+sumram[11][129]+sumram[11][130]+sumram[11][131]+sumram[11][132]+sumram[11][133]+sumram[11][134]+sumram[11][135]+sumram[11][136];
    assign sumcache[12]=sumram[12][0]+sumram[12][1]+sumram[12][2]+sumram[12][3]+sumram[12][4]+sumram[12][5]+sumram[12][6]+sumram[12][7]+sumram[12][8]+sumram[12][9]+sumram[12][10]+sumram[12][11]+sumram[12][12]+sumram[12][13]+sumram[12][14]+sumram[12][15]+sumram[12][16]+sumram[12][17]+sumram[12][18]+sumram[12][19]+sumram[12][20]+sumram[12][21]+sumram[12][22]+sumram[12][23]+sumram[12][24]+sumram[12][25]+sumram[12][26]+sumram[12][27]+sumram[12][28]+sumram[12][29]+sumram[12][30]+sumram[12][31]+sumram[12][32]+sumram[12][33]+sumram[12][34]+sumram[12][35]+sumram[12][36]+sumram[12][37]+sumram[12][38]+sumram[12][39]+sumram[12][40]+sumram[12][41]+sumram[12][42]+sumram[12][43]+sumram[12][44]+sumram[12][45]+sumram[12][46]+sumram[12][47]+sumram[12][48]+sumram[12][49]+sumram[12][50]+sumram[12][51]+sumram[12][52]+sumram[12][53]+sumram[12][54]+sumram[12][55]+sumram[12][56]+sumram[12][57]+sumram[12][58]+sumram[12][59]+sumram[12][60]+sumram[12][61]+sumram[12][62]+sumram[12][63]+sumram[12][64]+sumram[12][65]+sumram[12][66]+sumram[12][67]+sumram[12][68]+sumram[12][69]+sumram[12][70]+sumram[12][71]+sumram[12][72]+sumram[12][73]+sumram[12][74]+sumram[12][75]+sumram[12][76]+sumram[12][77]+sumram[12][78]+sumram[12][79]+sumram[12][80]+sumram[12][81]+sumram[12][82]+sumram[12][83]+sumram[12][84]+sumram[12][85]+sumram[12][86]+sumram[12][87]+sumram[12][88]+sumram[12][89]+sumram[12][90]+sumram[12][91]+sumram[12][92]+sumram[12][93]+sumram[12][94]+sumram[12][95]+sumram[12][96]+sumram[12][97]+sumram[12][98]+sumram[12][99]+sumram[12][100]+sumram[12][101]+sumram[12][102]+sumram[12][103]+sumram[12][104]+sumram[12][105]+sumram[12][106]+sumram[12][107]+sumram[12][108]+sumram[12][109]+sumram[12][110]+sumram[12][111]+sumram[12][112]+sumram[12][113]+sumram[12][114]+sumram[12][115]+sumram[12][116]+sumram[12][117]+sumram[12][118]+sumram[12][119]+sumram[12][120]+sumram[12][121]+sumram[12][122]+sumram[12][123]+sumram[12][124]+sumram[12][125]+sumram[12][126]+sumram[12][127]+sumram[12][128]+sumram[12][129]+sumram[12][130]+sumram[12][131]+sumram[12][132]+sumram[12][133]+sumram[12][134]+sumram[12][135]+sumram[12][136];
    assign sumcache[13]=sumram[13][0]+sumram[13][1]+sumram[13][2]+sumram[13][3]+sumram[13][4]+sumram[13][5]+sumram[13][6]+sumram[13][7]+sumram[13][8]+sumram[13][9]+sumram[13][10]+sumram[13][11]+sumram[13][12]+sumram[13][13]+sumram[13][14]+sumram[13][15]+sumram[13][16]+sumram[13][17]+sumram[13][18]+sumram[13][19]+sumram[13][20]+sumram[13][21]+sumram[13][22]+sumram[13][23]+sumram[13][24]+sumram[13][25]+sumram[13][26]+sumram[13][27]+sumram[13][28]+sumram[13][29]+sumram[13][30]+sumram[13][31]+sumram[13][32]+sumram[13][33]+sumram[13][34]+sumram[13][35]+sumram[13][36]+sumram[13][37]+sumram[13][38]+sumram[13][39]+sumram[13][40]+sumram[13][41]+sumram[13][42]+sumram[13][43]+sumram[13][44]+sumram[13][45]+sumram[13][46]+sumram[13][47]+sumram[13][48]+sumram[13][49]+sumram[13][50]+sumram[13][51]+sumram[13][52]+sumram[13][53]+sumram[13][54]+sumram[13][55]+sumram[13][56]+sumram[13][57]+sumram[13][58]+sumram[13][59]+sumram[13][60]+sumram[13][61]+sumram[13][62]+sumram[13][63]+sumram[13][64]+sumram[13][65]+sumram[13][66]+sumram[13][67]+sumram[13][68]+sumram[13][69]+sumram[13][70]+sumram[13][71]+sumram[13][72]+sumram[13][73]+sumram[13][74]+sumram[13][75]+sumram[13][76]+sumram[13][77]+sumram[13][78]+sumram[13][79]+sumram[13][80]+sumram[13][81]+sumram[13][82]+sumram[13][83]+sumram[13][84]+sumram[13][85]+sumram[13][86]+sumram[13][87]+sumram[13][88]+sumram[13][89]+sumram[13][90]+sumram[13][91]+sumram[13][92]+sumram[13][93]+sumram[13][94]+sumram[13][95]+sumram[13][96]+sumram[13][97]+sumram[13][98]+sumram[13][99]+sumram[13][100]+sumram[13][101]+sumram[13][102]+sumram[13][103]+sumram[13][104]+sumram[13][105]+sumram[13][106]+sumram[13][107]+sumram[13][108]+sumram[13][109]+sumram[13][110]+sumram[13][111]+sumram[13][112]+sumram[13][113]+sumram[13][114]+sumram[13][115]+sumram[13][116]+sumram[13][117]+sumram[13][118]+sumram[13][119]+sumram[13][120]+sumram[13][121]+sumram[13][122]+sumram[13][123]+sumram[13][124]+sumram[13][125]+sumram[13][126]+sumram[13][127]+sumram[13][128]+sumram[13][129]+sumram[13][130]+sumram[13][131]+sumram[13][132]+sumram[13][133]+sumram[13][134]+sumram[13][135]+sumram[13][136];
    assign sumcache[14]=sumram[14][0]+sumram[14][1]+sumram[14][2]+sumram[14][3]+sumram[14][4]+sumram[14][5]+sumram[14][6]+sumram[14][7]+sumram[14][8]+sumram[14][9]+sumram[14][10]+sumram[14][11]+sumram[14][12]+sumram[14][13]+sumram[14][14]+sumram[14][15]+sumram[14][16]+sumram[14][17]+sumram[14][18]+sumram[14][19]+sumram[14][20]+sumram[14][21]+sumram[14][22]+sumram[14][23]+sumram[14][24]+sumram[14][25]+sumram[14][26]+sumram[14][27]+sumram[14][28]+sumram[14][29]+sumram[14][30]+sumram[14][31]+sumram[14][32]+sumram[14][33]+sumram[14][34]+sumram[14][35]+sumram[14][36]+sumram[14][37]+sumram[14][38]+sumram[14][39]+sumram[14][40]+sumram[14][41]+sumram[14][42]+sumram[14][43]+sumram[14][44]+sumram[14][45]+sumram[14][46]+sumram[14][47]+sumram[14][48]+sumram[14][49]+sumram[14][50]+sumram[14][51]+sumram[14][52]+sumram[14][53]+sumram[14][54]+sumram[14][55]+sumram[14][56]+sumram[14][57]+sumram[14][58]+sumram[14][59]+sumram[14][60]+sumram[14][61]+sumram[14][62]+sumram[14][63]+sumram[14][64]+sumram[14][65]+sumram[14][66]+sumram[14][67]+sumram[14][68]+sumram[14][69]+sumram[14][70]+sumram[14][71]+sumram[14][72]+sumram[14][73]+sumram[14][74]+sumram[14][75]+sumram[14][76]+sumram[14][77]+sumram[14][78]+sumram[14][79]+sumram[14][80]+sumram[14][81]+sumram[14][82]+sumram[14][83]+sumram[14][84]+sumram[14][85]+sumram[14][86]+sumram[14][87]+sumram[14][88]+sumram[14][89]+sumram[14][90]+sumram[14][91]+sumram[14][92]+sumram[14][93]+sumram[14][94]+sumram[14][95]+sumram[14][96]+sumram[14][97]+sumram[14][98]+sumram[14][99]+sumram[14][100]+sumram[14][101]+sumram[14][102]+sumram[14][103]+sumram[14][104]+sumram[14][105]+sumram[14][106]+sumram[14][107]+sumram[14][108]+sumram[14][109]+sumram[14][110]+sumram[14][111]+sumram[14][112]+sumram[14][113]+sumram[14][114]+sumram[14][115]+sumram[14][116]+sumram[14][117]+sumram[14][118]+sumram[14][119]+sumram[14][120]+sumram[14][121]+sumram[14][122]+sumram[14][123]+sumram[14][124]+sumram[14][125]+sumram[14][126]+sumram[14][127]+sumram[14][128]+sumram[14][129]+sumram[14][130]+sumram[14][131]+sumram[14][132]+sumram[14][133]+sumram[14][134]+sumram[14][135]+sumram[14][136];
    assign sumcache[15]=sumram[15][0]+sumram[15][1]+sumram[15][2]+sumram[15][3]+sumram[15][4]+sumram[15][5]+sumram[15][6]+sumram[15][7]+sumram[15][8]+sumram[15][9]+sumram[15][10]+sumram[15][11]+sumram[15][12]+sumram[15][13]+sumram[15][14]+sumram[15][15]+sumram[15][16]+sumram[15][17]+sumram[15][18]+sumram[15][19]+sumram[15][20]+sumram[15][21]+sumram[15][22]+sumram[15][23]+sumram[15][24]+sumram[15][25]+sumram[15][26]+sumram[15][27]+sumram[15][28]+sumram[15][29]+sumram[15][30]+sumram[15][31]+sumram[15][32]+sumram[15][33]+sumram[15][34]+sumram[15][35]+sumram[15][36]+sumram[15][37]+sumram[15][38]+sumram[15][39]+sumram[15][40]+sumram[15][41]+sumram[15][42]+sumram[15][43]+sumram[15][44]+sumram[15][45]+sumram[15][46]+sumram[15][47]+sumram[15][48]+sumram[15][49]+sumram[15][50]+sumram[15][51]+sumram[15][52]+sumram[15][53]+sumram[15][54]+sumram[15][55]+sumram[15][56]+sumram[15][57]+sumram[15][58]+sumram[15][59]+sumram[15][60]+sumram[15][61]+sumram[15][62]+sumram[15][63]+sumram[15][64]+sumram[15][65]+sumram[15][66]+sumram[15][67]+sumram[15][68]+sumram[15][69]+sumram[15][70]+sumram[15][71]+sumram[15][72]+sumram[15][73]+sumram[15][74]+sumram[15][75]+sumram[15][76]+sumram[15][77]+sumram[15][78]+sumram[15][79]+sumram[15][80]+sumram[15][81]+sumram[15][82]+sumram[15][83]+sumram[15][84]+sumram[15][85]+sumram[15][86]+sumram[15][87]+sumram[15][88]+sumram[15][89]+sumram[15][90]+sumram[15][91]+sumram[15][92]+sumram[15][93]+sumram[15][94]+sumram[15][95]+sumram[15][96]+sumram[15][97]+sumram[15][98]+sumram[15][99]+sumram[15][100]+sumram[15][101]+sumram[15][102]+sumram[15][103]+sumram[15][104]+sumram[15][105]+sumram[15][106]+sumram[15][107]+sumram[15][108]+sumram[15][109]+sumram[15][110]+sumram[15][111]+sumram[15][112]+sumram[15][113]+sumram[15][114]+sumram[15][115]+sumram[15][116]+sumram[15][117]+sumram[15][118]+sumram[15][119]+sumram[15][120]+sumram[15][121]+sumram[15][122]+sumram[15][123]+sumram[15][124]+sumram[15][125]+sumram[15][126]+sumram[15][127]+sumram[15][128]+sumram[15][129]+sumram[15][130]+sumram[15][131]+sumram[15][132]+sumram[15][133]+sumram[15][134]+sumram[15][135]+sumram[15][136];
    assign sumcache[16]=sumram[16][0]+sumram[16][1]+sumram[16][2]+sumram[16][3]+sumram[16][4]+sumram[16][5]+sumram[16][6]+sumram[16][7]+sumram[16][8]+sumram[16][9]+sumram[16][10]+sumram[16][11]+sumram[16][12]+sumram[16][13]+sumram[16][14]+sumram[16][15]+sumram[16][16]+sumram[16][17]+sumram[16][18]+sumram[16][19]+sumram[16][20]+sumram[16][21]+sumram[16][22]+sumram[16][23]+sumram[16][24]+sumram[16][25]+sumram[16][26]+sumram[16][27]+sumram[16][28]+sumram[16][29]+sumram[16][30]+sumram[16][31]+sumram[16][32]+sumram[16][33]+sumram[16][34]+sumram[16][35]+sumram[16][36]+sumram[16][37]+sumram[16][38]+sumram[16][39]+sumram[16][40]+sumram[16][41]+sumram[16][42]+sumram[16][43]+sumram[16][44]+sumram[16][45]+sumram[16][46]+sumram[16][47]+sumram[16][48]+sumram[16][49]+sumram[16][50]+sumram[16][51]+sumram[16][52]+sumram[16][53]+sumram[16][54]+sumram[16][55]+sumram[16][56]+sumram[16][57]+sumram[16][58]+sumram[16][59]+sumram[16][60]+sumram[16][61]+sumram[16][62]+sumram[16][63]+sumram[16][64]+sumram[16][65]+sumram[16][66]+sumram[16][67]+sumram[16][68]+sumram[16][69]+sumram[16][70]+sumram[16][71]+sumram[16][72]+sumram[16][73]+sumram[16][74]+sumram[16][75]+sumram[16][76]+sumram[16][77]+sumram[16][78]+sumram[16][79]+sumram[16][80]+sumram[16][81]+sumram[16][82]+sumram[16][83]+sumram[16][84]+sumram[16][85]+sumram[16][86]+sumram[16][87]+sumram[16][88]+sumram[16][89]+sumram[16][90]+sumram[16][91]+sumram[16][92]+sumram[16][93]+sumram[16][94]+sumram[16][95]+sumram[16][96]+sumram[16][97]+sumram[16][98]+sumram[16][99]+sumram[16][100]+sumram[16][101]+sumram[16][102]+sumram[16][103]+sumram[16][104]+sumram[16][105]+sumram[16][106]+sumram[16][107]+sumram[16][108]+sumram[16][109]+sumram[16][110]+sumram[16][111]+sumram[16][112]+sumram[16][113]+sumram[16][114]+sumram[16][115]+sumram[16][116]+sumram[16][117]+sumram[16][118]+sumram[16][119]+sumram[16][120]+sumram[16][121]+sumram[16][122]+sumram[16][123]+sumram[16][124]+sumram[16][125]+sumram[16][126]+sumram[16][127]+sumram[16][128]+sumram[16][129]+sumram[16][130]+sumram[16][131]+sumram[16][132]+sumram[16][133]+sumram[16][134]+sumram[16][135]+sumram[16][136];
    assign sumcache[17]=sumram[17][0]+sumram[17][1]+sumram[17][2]+sumram[17][3]+sumram[17][4]+sumram[17][5]+sumram[17][6]+sumram[17][7]+sumram[17][8]+sumram[17][9]+sumram[17][10]+sumram[17][11]+sumram[17][12]+sumram[17][13]+sumram[17][14]+sumram[17][15]+sumram[17][16]+sumram[17][17]+sumram[17][18]+sumram[17][19]+sumram[17][20]+sumram[17][21]+sumram[17][22]+sumram[17][23]+sumram[17][24]+sumram[17][25]+sumram[17][26]+sumram[17][27]+sumram[17][28]+sumram[17][29]+sumram[17][30]+sumram[17][31]+sumram[17][32]+sumram[17][33]+sumram[17][34]+sumram[17][35]+sumram[17][36]+sumram[17][37]+sumram[17][38]+sumram[17][39]+sumram[17][40]+sumram[17][41]+sumram[17][42]+sumram[17][43]+sumram[17][44]+sumram[17][45]+sumram[17][46]+sumram[17][47]+sumram[17][48]+sumram[17][49]+sumram[17][50]+sumram[17][51]+sumram[17][52]+sumram[17][53]+sumram[17][54]+sumram[17][55]+sumram[17][56]+sumram[17][57]+sumram[17][58]+sumram[17][59]+sumram[17][60]+sumram[17][61]+sumram[17][62]+sumram[17][63]+sumram[17][64]+sumram[17][65]+sumram[17][66]+sumram[17][67]+sumram[17][68]+sumram[17][69]+sumram[17][70]+sumram[17][71]+sumram[17][72]+sumram[17][73]+sumram[17][74]+sumram[17][75]+sumram[17][76]+sumram[17][77]+sumram[17][78]+sumram[17][79]+sumram[17][80]+sumram[17][81]+sumram[17][82]+sumram[17][83]+sumram[17][84]+sumram[17][85]+sumram[17][86]+sumram[17][87]+sumram[17][88]+sumram[17][89]+sumram[17][90]+sumram[17][91]+sumram[17][92]+sumram[17][93]+sumram[17][94]+sumram[17][95]+sumram[17][96]+sumram[17][97]+sumram[17][98]+sumram[17][99]+sumram[17][100]+sumram[17][101]+sumram[17][102]+sumram[17][103]+sumram[17][104]+sumram[17][105]+sumram[17][106]+sumram[17][107]+sumram[17][108]+sumram[17][109]+sumram[17][110]+sumram[17][111]+sumram[17][112]+sumram[17][113]+sumram[17][114]+sumram[17][115]+sumram[17][116]+sumram[17][117]+sumram[17][118]+sumram[17][119]+sumram[17][120]+sumram[17][121]+sumram[17][122]+sumram[17][123]+sumram[17][124]+sumram[17][125]+sumram[17][126]+sumram[17][127]+sumram[17][128]+sumram[17][129]+sumram[17][130]+sumram[17][131]+sumram[17][132]+sumram[17][133]+sumram[17][134]+sumram[17][135]+sumram[17][136];
    assign sumcache[18]=sumram[18][0]+sumram[18][1]+sumram[18][2]+sumram[18][3]+sumram[18][4]+sumram[18][5]+sumram[18][6]+sumram[18][7]+sumram[18][8]+sumram[18][9]+sumram[18][10]+sumram[18][11]+sumram[18][12]+sumram[18][13]+sumram[18][14]+sumram[18][15]+sumram[18][16]+sumram[18][17]+sumram[18][18]+sumram[18][19]+sumram[18][20]+sumram[18][21]+sumram[18][22]+sumram[18][23]+sumram[18][24]+sumram[18][25]+sumram[18][26]+sumram[18][27]+sumram[18][28]+sumram[18][29]+sumram[18][30]+sumram[18][31]+sumram[18][32]+sumram[18][33]+sumram[18][34]+sumram[18][35]+sumram[18][36]+sumram[18][37]+sumram[18][38]+sumram[18][39]+sumram[18][40]+sumram[18][41]+sumram[18][42]+sumram[18][43]+sumram[18][44]+sumram[18][45]+sumram[18][46]+sumram[18][47]+sumram[18][48]+sumram[18][49]+sumram[18][50]+sumram[18][51]+sumram[18][52]+sumram[18][53]+sumram[18][54]+sumram[18][55]+sumram[18][56]+sumram[18][57]+sumram[18][58]+sumram[18][59]+sumram[18][60]+sumram[18][61]+sumram[18][62]+sumram[18][63]+sumram[18][64]+sumram[18][65]+sumram[18][66]+sumram[18][67]+sumram[18][68]+sumram[18][69]+sumram[18][70]+sumram[18][71]+sumram[18][72]+sumram[18][73]+sumram[18][74]+sumram[18][75]+sumram[18][76]+sumram[18][77]+sumram[18][78]+sumram[18][79]+sumram[18][80]+sumram[18][81]+sumram[18][82]+sumram[18][83]+sumram[18][84]+sumram[18][85]+sumram[18][86]+sumram[18][87]+sumram[18][88]+sumram[18][89]+sumram[18][90]+sumram[18][91]+sumram[18][92]+sumram[18][93]+sumram[18][94]+sumram[18][95]+sumram[18][96]+sumram[18][97]+sumram[18][98]+sumram[18][99]+sumram[18][100]+sumram[18][101]+sumram[18][102]+sumram[18][103]+sumram[18][104]+sumram[18][105]+sumram[18][106]+sumram[18][107]+sumram[18][108]+sumram[18][109]+sumram[18][110]+sumram[18][111]+sumram[18][112]+sumram[18][113]+sumram[18][114]+sumram[18][115]+sumram[18][116]+sumram[18][117]+sumram[18][118]+sumram[18][119]+sumram[18][120]+sumram[18][121]+sumram[18][122]+sumram[18][123]+sumram[18][124]+sumram[18][125]+sumram[18][126]+sumram[18][127]+sumram[18][128]+sumram[18][129]+sumram[18][130]+sumram[18][131]+sumram[18][132]+sumram[18][133]+sumram[18][134]+sumram[18][135]+sumram[18][136];
    assign sumcache[19]=sumram[19][0]+sumram[19][1]+sumram[19][2]+sumram[19][3]+sumram[19][4]+sumram[19][5]+sumram[19][6]+sumram[19][7]+sumram[19][8]+sumram[19][9]+sumram[19][10]+sumram[19][11]+sumram[19][12]+sumram[19][13]+sumram[19][14]+sumram[19][15]+sumram[19][16]+sumram[19][17]+sumram[19][18]+sumram[19][19]+sumram[19][20]+sumram[19][21]+sumram[19][22]+sumram[19][23]+sumram[19][24]+sumram[19][25]+sumram[19][26]+sumram[19][27]+sumram[19][28]+sumram[19][29]+sumram[19][30]+sumram[19][31]+sumram[19][32]+sumram[19][33]+sumram[19][34]+sumram[19][35]+sumram[19][36]+sumram[19][37]+sumram[19][38]+sumram[19][39]+sumram[19][40]+sumram[19][41]+sumram[19][42]+sumram[19][43]+sumram[19][44]+sumram[19][45]+sumram[19][46]+sumram[19][47]+sumram[19][48]+sumram[19][49]+sumram[19][50]+sumram[19][51]+sumram[19][52]+sumram[19][53]+sumram[19][54]+sumram[19][55]+sumram[19][56]+sumram[19][57]+sumram[19][58]+sumram[19][59]+sumram[19][60]+sumram[19][61]+sumram[19][62]+sumram[19][63]+sumram[19][64]+sumram[19][65]+sumram[19][66]+sumram[19][67]+sumram[19][68]+sumram[19][69]+sumram[19][70]+sumram[19][71]+sumram[19][72]+sumram[19][73]+sumram[19][74]+sumram[19][75]+sumram[19][76]+sumram[19][77]+sumram[19][78]+sumram[19][79]+sumram[19][80]+sumram[19][81]+sumram[19][82]+sumram[19][83]+sumram[19][84]+sumram[19][85]+sumram[19][86]+sumram[19][87]+sumram[19][88]+sumram[19][89]+sumram[19][90]+sumram[19][91]+sumram[19][92]+sumram[19][93]+sumram[19][94]+sumram[19][95]+sumram[19][96]+sumram[19][97]+sumram[19][98]+sumram[19][99]+sumram[19][100]+sumram[19][101]+sumram[19][102]+sumram[19][103]+sumram[19][104]+sumram[19][105]+sumram[19][106]+sumram[19][107]+sumram[19][108]+sumram[19][109]+sumram[19][110]+sumram[19][111]+sumram[19][112]+sumram[19][113]+sumram[19][114]+sumram[19][115]+sumram[19][116]+sumram[19][117]+sumram[19][118]+sumram[19][119]+sumram[19][120]+sumram[19][121]+sumram[19][122]+sumram[19][123]+sumram[19][124]+sumram[19][125]+sumram[19][126]+sumram[19][127]+sumram[19][128]+sumram[19][129]+sumram[19][130]+sumram[19][131]+sumram[19][132]+sumram[19][133]+sumram[19][134]+sumram[19][135]+sumram[19][136];
    assign sumcache[20]=sumram[20][0]+sumram[20][1]+sumram[20][2]+sumram[20][3]+sumram[20][4]+sumram[20][5]+sumram[20][6]+sumram[20][7]+sumram[20][8]+sumram[20][9]+sumram[20][10]+sumram[20][11]+sumram[20][12]+sumram[20][13]+sumram[20][14]+sumram[20][15]+sumram[20][16]+sumram[20][17]+sumram[20][18]+sumram[20][19]+sumram[20][20]+sumram[20][21]+sumram[20][22]+sumram[20][23]+sumram[20][24]+sumram[20][25]+sumram[20][26]+sumram[20][27]+sumram[20][28]+sumram[20][29]+sumram[20][30]+sumram[20][31]+sumram[20][32]+sumram[20][33]+sumram[20][34]+sumram[20][35]+sumram[20][36]+sumram[20][37]+sumram[20][38]+sumram[20][39]+sumram[20][40]+sumram[20][41]+sumram[20][42]+sumram[20][43]+sumram[20][44]+sumram[20][45]+sumram[20][46]+sumram[20][47]+sumram[20][48]+sumram[20][49]+sumram[20][50]+sumram[20][51]+sumram[20][52]+sumram[20][53]+sumram[20][54]+sumram[20][55]+sumram[20][56]+sumram[20][57]+sumram[20][58]+sumram[20][59]+sumram[20][60]+sumram[20][61]+sumram[20][62]+sumram[20][63]+sumram[20][64]+sumram[20][65]+sumram[20][66]+sumram[20][67]+sumram[20][68]+sumram[20][69]+sumram[20][70]+sumram[20][71]+sumram[20][72]+sumram[20][73]+sumram[20][74]+sumram[20][75]+sumram[20][76]+sumram[20][77]+sumram[20][78]+sumram[20][79]+sumram[20][80]+sumram[20][81]+sumram[20][82]+sumram[20][83]+sumram[20][84]+sumram[20][85]+sumram[20][86]+sumram[20][87]+sumram[20][88]+sumram[20][89]+sumram[20][90]+sumram[20][91]+sumram[20][92]+sumram[20][93]+sumram[20][94]+sumram[20][95]+sumram[20][96]+sumram[20][97]+sumram[20][98]+sumram[20][99]+sumram[20][100]+sumram[20][101]+sumram[20][102]+sumram[20][103]+sumram[20][104]+sumram[20][105]+sumram[20][106]+sumram[20][107]+sumram[20][108]+sumram[20][109]+sumram[20][110]+sumram[20][111]+sumram[20][112]+sumram[20][113]+sumram[20][114]+sumram[20][115]+sumram[20][116]+sumram[20][117]+sumram[20][118]+sumram[20][119]+sumram[20][120]+sumram[20][121]+sumram[20][122]+sumram[20][123]+sumram[20][124]+sumram[20][125]+sumram[20][126]+sumram[20][127]+sumram[20][128]+sumram[20][129]+sumram[20][130]+sumram[20][131]+sumram[20][132]+sumram[20][133]+sumram[20][134]+sumram[20][135]+sumram[20][136];
    assign sumcache[21]=sumram[21][0]+sumram[21][1]+sumram[21][2]+sumram[21][3]+sumram[21][4]+sumram[21][5]+sumram[21][6]+sumram[21][7]+sumram[21][8]+sumram[21][9]+sumram[21][10]+sumram[21][11]+sumram[21][12]+sumram[21][13]+sumram[21][14]+sumram[21][15]+sumram[21][16]+sumram[21][17]+sumram[21][18]+sumram[21][19]+sumram[21][20]+sumram[21][21]+sumram[21][22]+sumram[21][23]+sumram[21][24]+sumram[21][25]+sumram[21][26]+sumram[21][27]+sumram[21][28]+sumram[21][29]+sumram[21][30]+sumram[21][31]+sumram[21][32]+sumram[21][33]+sumram[21][34]+sumram[21][35]+sumram[21][36]+sumram[21][37]+sumram[21][38]+sumram[21][39]+sumram[21][40]+sumram[21][41]+sumram[21][42]+sumram[21][43]+sumram[21][44]+sumram[21][45]+sumram[21][46]+sumram[21][47]+sumram[21][48]+sumram[21][49]+sumram[21][50]+sumram[21][51]+sumram[21][52]+sumram[21][53]+sumram[21][54]+sumram[21][55]+sumram[21][56]+sumram[21][57]+sumram[21][58]+sumram[21][59]+sumram[21][60]+sumram[21][61]+sumram[21][62]+sumram[21][63]+sumram[21][64]+sumram[21][65]+sumram[21][66]+sumram[21][67]+sumram[21][68]+sumram[21][69]+sumram[21][70]+sumram[21][71]+sumram[21][72]+sumram[21][73]+sumram[21][74]+sumram[21][75]+sumram[21][76]+sumram[21][77]+sumram[21][78]+sumram[21][79]+sumram[21][80]+sumram[21][81]+sumram[21][82]+sumram[21][83]+sumram[21][84]+sumram[21][85]+sumram[21][86]+sumram[21][87]+sumram[21][88]+sumram[21][89]+sumram[21][90]+sumram[21][91]+sumram[21][92]+sumram[21][93]+sumram[21][94]+sumram[21][95]+sumram[21][96]+sumram[21][97]+sumram[21][98]+sumram[21][99]+sumram[21][100]+sumram[21][101]+sumram[21][102]+sumram[21][103]+sumram[21][104]+sumram[21][105]+sumram[21][106]+sumram[21][107]+sumram[21][108]+sumram[21][109]+sumram[21][110]+sumram[21][111]+sumram[21][112]+sumram[21][113]+sumram[21][114]+sumram[21][115]+sumram[21][116]+sumram[21][117]+sumram[21][118]+sumram[21][119]+sumram[21][120]+sumram[21][121]+sumram[21][122]+sumram[21][123]+sumram[21][124]+sumram[21][125]+sumram[21][126]+sumram[21][127]+sumram[21][128]+sumram[21][129]+sumram[21][130]+sumram[21][131]+sumram[21][132]+sumram[21][133]+sumram[21][134]+sumram[21][135]+sumram[21][136];
    assign sumcache[22]=sumram[22][0]+sumram[22][1]+sumram[22][2]+sumram[22][3]+sumram[22][4]+sumram[22][5]+sumram[22][6]+sumram[22][7]+sumram[22][8]+sumram[22][9]+sumram[22][10]+sumram[22][11]+sumram[22][12]+sumram[22][13]+sumram[22][14]+sumram[22][15]+sumram[22][16]+sumram[22][17]+sumram[22][18]+sumram[22][19]+sumram[22][20]+sumram[22][21]+sumram[22][22]+sumram[22][23]+sumram[22][24]+sumram[22][25]+sumram[22][26]+sumram[22][27]+sumram[22][28]+sumram[22][29]+sumram[22][30]+sumram[22][31]+sumram[22][32]+sumram[22][33]+sumram[22][34]+sumram[22][35]+sumram[22][36]+sumram[22][37]+sumram[22][38]+sumram[22][39]+sumram[22][40]+sumram[22][41]+sumram[22][42]+sumram[22][43]+sumram[22][44]+sumram[22][45]+sumram[22][46]+sumram[22][47]+sumram[22][48]+sumram[22][49]+sumram[22][50]+sumram[22][51]+sumram[22][52]+sumram[22][53]+sumram[22][54]+sumram[22][55]+sumram[22][56]+sumram[22][57]+sumram[22][58]+sumram[22][59]+sumram[22][60]+sumram[22][61]+sumram[22][62]+sumram[22][63]+sumram[22][64]+sumram[22][65]+sumram[22][66]+sumram[22][67]+sumram[22][68]+sumram[22][69]+sumram[22][70]+sumram[22][71]+sumram[22][72]+sumram[22][73]+sumram[22][74]+sumram[22][75]+sumram[22][76]+sumram[22][77]+sumram[22][78]+sumram[22][79]+sumram[22][80]+sumram[22][81]+sumram[22][82]+sumram[22][83]+sumram[22][84]+sumram[22][85]+sumram[22][86]+sumram[22][87]+sumram[22][88]+sumram[22][89]+sumram[22][90]+sumram[22][91]+sumram[22][92]+sumram[22][93]+sumram[22][94]+sumram[22][95]+sumram[22][96]+sumram[22][97]+sumram[22][98]+sumram[22][99]+sumram[22][100]+sumram[22][101]+sumram[22][102]+sumram[22][103]+sumram[22][104]+sumram[22][105]+sumram[22][106]+sumram[22][107]+sumram[22][108]+sumram[22][109]+sumram[22][110]+sumram[22][111]+sumram[22][112]+sumram[22][113]+sumram[22][114]+sumram[22][115]+sumram[22][116]+sumram[22][117]+sumram[22][118]+sumram[22][119]+sumram[22][120]+sumram[22][121]+sumram[22][122]+sumram[22][123]+sumram[22][124]+sumram[22][125]+sumram[22][126]+sumram[22][127]+sumram[22][128]+sumram[22][129]+sumram[22][130]+sumram[22][131]+sumram[22][132]+sumram[22][133]+sumram[22][134]+sumram[22][135]+sumram[22][136];
    assign sumcache[23]=sumram[23][0]+sumram[23][1]+sumram[23][2]+sumram[23][3]+sumram[23][4]+sumram[23][5]+sumram[23][6]+sumram[23][7]+sumram[23][8]+sumram[23][9]+sumram[23][10]+sumram[23][11]+sumram[23][12]+sumram[23][13]+sumram[23][14]+sumram[23][15]+sumram[23][16]+sumram[23][17]+sumram[23][18]+sumram[23][19]+sumram[23][20]+sumram[23][21]+sumram[23][22]+sumram[23][23]+sumram[23][24]+sumram[23][25]+sumram[23][26]+sumram[23][27]+sumram[23][28]+sumram[23][29]+sumram[23][30]+sumram[23][31]+sumram[23][32]+sumram[23][33]+sumram[23][34]+sumram[23][35]+sumram[23][36]+sumram[23][37]+sumram[23][38]+sumram[23][39]+sumram[23][40]+sumram[23][41]+sumram[23][42]+sumram[23][43]+sumram[23][44]+sumram[23][45]+sumram[23][46]+sumram[23][47]+sumram[23][48]+sumram[23][49]+sumram[23][50]+sumram[23][51]+sumram[23][52]+sumram[23][53]+sumram[23][54]+sumram[23][55]+sumram[23][56]+sumram[23][57]+sumram[23][58]+sumram[23][59]+sumram[23][60]+sumram[23][61]+sumram[23][62]+sumram[23][63]+sumram[23][64]+sumram[23][65]+sumram[23][66]+sumram[23][67]+sumram[23][68]+sumram[23][69]+sumram[23][70]+sumram[23][71]+sumram[23][72]+sumram[23][73]+sumram[23][74]+sumram[23][75]+sumram[23][76]+sumram[23][77]+sumram[23][78]+sumram[23][79]+sumram[23][80]+sumram[23][81]+sumram[23][82]+sumram[23][83]+sumram[23][84]+sumram[23][85]+sumram[23][86]+sumram[23][87]+sumram[23][88]+sumram[23][89]+sumram[23][90]+sumram[23][91]+sumram[23][92]+sumram[23][93]+sumram[23][94]+sumram[23][95]+sumram[23][96]+sumram[23][97]+sumram[23][98]+sumram[23][99]+sumram[23][100]+sumram[23][101]+sumram[23][102]+sumram[23][103]+sumram[23][104]+sumram[23][105]+sumram[23][106]+sumram[23][107]+sumram[23][108]+sumram[23][109]+sumram[23][110]+sumram[23][111]+sumram[23][112]+sumram[23][113]+sumram[23][114]+sumram[23][115]+sumram[23][116]+sumram[23][117]+sumram[23][118]+sumram[23][119]+sumram[23][120]+sumram[23][121]+sumram[23][122]+sumram[23][123]+sumram[23][124]+sumram[23][125]+sumram[23][126]+sumram[23][127]+sumram[23][128]+sumram[23][129]+sumram[23][130]+sumram[23][131]+sumram[23][132]+sumram[23][133]+sumram[23][134]+sumram[23][135]+sumram[23][136];
    assign sumcache[24]=sumram[24][0]+sumram[24][1]+sumram[24][2]+sumram[24][3]+sumram[24][4]+sumram[24][5]+sumram[24][6]+sumram[24][7]+sumram[24][8]+sumram[24][9]+sumram[24][10]+sumram[24][11]+sumram[24][12]+sumram[24][13]+sumram[24][14]+sumram[24][15]+sumram[24][16]+sumram[24][17]+sumram[24][18]+sumram[24][19]+sumram[24][20]+sumram[24][21]+sumram[24][22]+sumram[24][23]+sumram[24][24]+sumram[24][25]+sumram[24][26]+sumram[24][27]+sumram[24][28]+sumram[24][29]+sumram[24][30]+sumram[24][31]+sumram[24][32]+sumram[24][33]+sumram[24][34]+sumram[24][35]+sumram[24][36]+sumram[24][37]+sumram[24][38]+sumram[24][39]+sumram[24][40]+sumram[24][41]+sumram[24][42]+sumram[24][43]+sumram[24][44]+sumram[24][45]+sumram[24][46]+sumram[24][47]+sumram[24][48]+sumram[24][49]+sumram[24][50]+sumram[24][51]+sumram[24][52]+sumram[24][53]+sumram[24][54]+sumram[24][55]+sumram[24][56]+sumram[24][57]+sumram[24][58]+sumram[24][59]+sumram[24][60]+sumram[24][61]+sumram[24][62]+sumram[24][63]+sumram[24][64]+sumram[24][65]+sumram[24][66]+sumram[24][67]+sumram[24][68]+sumram[24][69]+sumram[24][70]+sumram[24][71]+sumram[24][72]+sumram[24][73]+sumram[24][74]+sumram[24][75]+sumram[24][76]+sumram[24][77]+sumram[24][78]+sumram[24][79]+sumram[24][80]+sumram[24][81]+sumram[24][82]+sumram[24][83]+sumram[24][84]+sumram[24][85]+sumram[24][86]+sumram[24][87]+sumram[24][88]+sumram[24][89]+sumram[24][90]+sumram[24][91]+sumram[24][92]+sumram[24][93]+sumram[24][94]+sumram[24][95]+sumram[24][96]+sumram[24][97]+sumram[24][98]+sumram[24][99]+sumram[24][100]+sumram[24][101]+sumram[24][102]+sumram[24][103]+sumram[24][104]+sumram[24][105]+sumram[24][106]+sumram[24][107]+sumram[24][108]+sumram[24][109]+sumram[24][110]+sumram[24][111]+sumram[24][112]+sumram[24][113]+sumram[24][114]+sumram[24][115]+sumram[24][116]+sumram[24][117]+sumram[24][118]+sumram[24][119]+sumram[24][120]+sumram[24][121]+sumram[24][122]+sumram[24][123]+sumram[24][124]+sumram[24][125]+sumram[24][126]+sumram[24][127]+sumram[24][128]+sumram[24][129]+sumram[24][130]+sumram[24][131]+sumram[24][132]+sumram[24][133]+sumram[24][134]+sumram[24][135]+sumram[24][136];
    assign sumcache[25]=sumram[25][0]+sumram[25][1]+sumram[25][2]+sumram[25][3]+sumram[25][4]+sumram[25][5]+sumram[25][6]+sumram[25][7]+sumram[25][8]+sumram[25][9]+sumram[25][10]+sumram[25][11]+sumram[25][12]+sumram[25][13]+sumram[25][14]+sumram[25][15]+sumram[25][16]+sumram[25][17]+sumram[25][18]+sumram[25][19]+sumram[25][20]+sumram[25][21]+sumram[25][22]+sumram[25][23]+sumram[25][24]+sumram[25][25]+sumram[25][26]+sumram[25][27]+sumram[25][28]+sumram[25][29]+sumram[25][30]+sumram[25][31]+sumram[25][32]+sumram[25][33]+sumram[25][34]+sumram[25][35]+sumram[25][36]+sumram[25][37]+sumram[25][38]+sumram[25][39]+sumram[25][40]+sumram[25][41]+sumram[25][42]+sumram[25][43]+sumram[25][44]+sumram[25][45]+sumram[25][46]+sumram[25][47]+sumram[25][48]+sumram[25][49]+sumram[25][50]+sumram[25][51]+sumram[25][52]+sumram[25][53]+sumram[25][54]+sumram[25][55]+sumram[25][56]+sumram[25][57]+sumram[25][58]+sumram[25][59]+sumram[25][60]+sumram[25][61]+sumram[25][62]+sumram[25][63]+sumram[25][64]+sumram[25][65]+sumram[25][66]+sumram[25][67]+sumram[25][68]+sumram[25][69]+sumram[25][70]+sumram[25][71]+sumram[25][72]+sumram[25][73]+sumram[25][74]+sumram[25][75]+sumram[25][76]+sumram[25][77]+sumram[25][78]+sumram[25][79]+sumram[25][80]+sumram[25][81]+sumram[25][82]+sumram[25][83]+sumram[25][84]+sumram[25][85]+sumram[25][86]+sumram[25][87]+sumram[25][88]+sumram[25][89]+sumram[25][90]+sumram[25][91]+sumram[25][92]+sumram[25][93]+sumram[25][94]+sumram[25][95]+sumram[25][96]+sumram[25][97]+sumram[25][98]+sumram[25][99]+sumram[25][100]+sumram[25][101]+sumram[25][102]+sumram[25][103]+sumram[25][104]+sumram[25][105]+sumram[25][106]+sumram[25][107]+sumram[25][108]+sumram[25][109]+sumram[25][110]+sumram[25][111]+sumram[25][112]+sumram[25][113]+sumram[25][114]+sumram[25][115]+sumram[25][116]+sumram[25][117]+sumram[25][118]+sumram[25][119]+sumram[25][120]+sumram[25][121]+sumram[25][122]+sumram[25][123]+sumram[25][124]+sumram[25][125]+sumram[25][126]+sumram[25][127]+sumram[25][128]+sumram[25][129]+sumram[25][130]+sumram[25][131]+sumram[25][132]+sumram[25][133]+sumram[25][134]+sumram[25][135]+sumram[25][136];
    assign sumcache[26]=sumram[26][0]+sumram[26][1]+sumram[26][2]+sumram[26][3]+sumram[26][4]+sumram[26][5]+sumram[26][6]+sumram[26][7]+sumram[26][8]+sumram[26][9]+sumram[26][10]+sumram[26][11]+sumram[26][12]+sumram[26][13]+sumram[26][14]+sumram[26][15]+sumram[26][16]+sumram[26][17]+sumram[26][18]+sumram[26][19]+sumram[26][20]+sumram[26][21]+sumram[26][22]+sumram[26][23]+sumram[26][24]+sumram[26][25]+sumram[26][26]+sumram[26][27]+sumram[26][28]+sumram[26][29]+sumram[26][30]+sumram[26][31]+sumram[26][32]+sumram[26][33]+sumram[26][34]+sumram[26][35]+sumram[26][36]+sumram[26][37]+sumram[26][38]+sumram[26][39]+sumram[26][40]+sumram[26][41]+sumram[26][42]+sumram[26][43]+sumram[26][44]+sumram[26][45]+sumram[26][46]+sumram[26][47]+sumram[26][48]+sumram[26][49]+sumram[26][50]+sumram[26][51]+sumram[26][52]+sumram[26][53]+sumram[26][54]+sumram[26][55]+sumram[26][56]+sumram[26][57]+sumram[26][58]+sumram[26][59]+sumram[26][60]+sumram[26][61]+sumram[26][62]+sumram[26][63]+sumram[26][64]+sumram[26][65]+sumram[26][66]+sumram[26][67]+sumram[26][68]+sumram[26][69]+sumram[26][70]+sumram[26][71]+sumram[26][72]+sumram[26][73]+sumram[26][74]+sumram[26][75]+sumram[26][76]+sumram[26][77]+sumram[26][78]+sumram[26][79]+sumram[26][80]+sumram[26][81]+sumram[26][82]+sumram[26][83]+sumram[26][84]+sumram[26][85]+sumram[26][86]+sumram[26][87]+sumram[26][88]+sumram[26][89]+sumram[26][90]+sumram[26][91]+sumram[26][92]+sumram[26][93]+sumram[26][94]+sumram[26][95]+sumram[26][96]+sumram[26][97]+sumram[26][98]+sumram[26][99]+sumram[26][100]+sumram[26][101]+sumram[26][102]+sumram[26][103]+sumram[26][104]+sumram[26][105]+sumram[26][106]+sumram[26][107]+sumram[26][108]+sumram[26][109]+sumram[26][110]+sumram[26][111]+sumram[26][112]+sumram[26][113]+sumram[26][114]+sumram[26][115]+sumram[26][116]+sumram[26][117]+sumram[26][118]+sumram[26][119]+sumram[26][120]+sumram[26][121]+sumram[26][122]+sumram[26][123]+sumram[26][124]+sumram[26][125]+sumram[26][126]+sumram[26][127]+sumram[26][128]+sumram[26][129]+sumram[26][130]+sumram[26][131]+sumram[26][132]+sumram[26][133]+sumram[26][134]+sumram[26][135]+sumram[26][136];
    assign sumcache[27]=sumram[27][0]+sumram[27][1]+sumram[27][2]+sumram[27][3]+sumram[27][4]+sumram[27][5]+sumram[27][6]+sumram[27][7]+sumram[27][8]+sumram[27][9]+sumram[27][10]+sumram[27][11]+sumram[27][12]+sumram[27][13]+sumram[27][14]+sumram[27][15]+sumram[27][16]+sumram[27][17]+sumram[27][18]+sumram[27][19]+sumram[27][20]+sumram[27][21]+sumram[27][22]+sumram[27][23]+sumram[27][24]+sumram[27][25]+sumram[27][26]+sumram[27][27]+sumram[27][28]+sumram[27][29]+sumram[27][30]+sumram[27][31]+sumram[27][32]+sumram[27][33]+sumram[27][34]+sumram[27][35]+sumram[27][36]+sumram[27][37]+sumram[27][38]+sumram[27][39]+sumram[27][40]+sumram[27][41]+sumram[27][42]+sumram[27][43]+sumram[27][44]+sumram[27][45]+sumram[27][46]+sumram[27][47]+sumram[27][48]+sumram[27][49]+sumram[27][50]+sumram[27][51]+sumram[27][52]+sumram[27][53]+sumram[27][54]+sumram[27][55]+sumram[27][56]+sumram[27][57]+sumram[27][58]+sumram[27][59]+sumram[27][60]+sumram[27][61]+sumram[27][62]+sumram[27][63]+sumram[27][64]+sumram[27][65]+sumram[27][66]+sumram[27][67]+sumram[27][68]+sumram[27][69]+sumram[27][70]+sumram[27][71]+sumram[27][72]+sumram[27][73]+sumram[27][74]+sumram[27][75]+sumram[27][76]+sumram[27][77]+sumram[27][78]+sumram[27][79]+sumram[27][80]+sumram[27][81]+sumram[27][82]+sumram[27][83]+sumram[27][84]+sumram[27][85]+sumram[27][86]+sumram[27][87]+sumram[27][88]+sumram[27][89]+sumram[27][90]+sumram[27][91]+sumram[27][92]+sumram[27][93]+sumram[27][94]+sumram[27][95]+sumram[27][96]+sumram[27][97]+sumram[27][98]+sumram[27][99]+sumram[27][100]+sumram[27][101]+sumram[27][102]+sumram[27][103]+sumram[27][104]+sumram[27][105]+sumram[27][106]+sumram[27][107]+sumram[27][108]+sumram[27][109]+sumram[27][110]+sumram[27][111]+sumram[27][112]+sumram[27][113]+sumram[27][114]+sumram[27][115]+sumram[27][116]+sumram[27][117]+sumram[27][118]+sumram[27][119]+sumram[27][120]+sumram[27][121]+sumram[27][122]+sumram[27][123]+sumram[27][124]+sumram[27][125]+sumram[27][126]+sumram[27][127]+sumram[27][128]+sumram[27][129]+sumram[27][130]+sumram[27][131]+sumram[27][132]+sumram[27][133]+sumram[27][134]+sumram[27][135]+sumram[27][136];
    assign sumcache[28]=sumram[28][0]+sumram[28][1]+sumram[28][2]+sumram[28][3]+sumram[28][4]+sumram[28][5]+sumram[28][6]+sumram[28][7]+sumram[28][8]+sumram[28][9]+sumram[28][10]+sumram[28][11]+sumram[28][12]+sumram[28][13]+sumram[28][14]+sumram[28][15]+sumram[28][16]+sumram[28][17]+sumram[28][18]+sumram[28][19]+sumram[28][20]+sumram[28][21]+sumram[28][22]+sumram[28][23]+sumram[28][24]+sumram[28][25]+sumram[28][26]+sumram[28][27]+sumram[28][28]+sumram[28][29]+sumram[28][30]+sumram[28][31]+sumram[28][32]+sumram[28][33]+sumram[28][34]+sumram[28][35]+sumram[28][36]+sumram[28][37]+sumram[28][38]+sumram[28][39]+sumram[28][40]+sumram[28][41]+sumram[28][42]+sumram[28][43]+sumram[28][44]+sumram[28][45]+sumram[28][46]+sumram[28][47]+sumram[28][48]+sumram[28][49]+sumram[28][50]+sumram[28][51]+sumram[28][52]+sumram[28][53]+sumram[28][54]+sumram[28][55]+sumram[28][56]+sumram[28][57]+sumram[28][58]+sumram[28][59]+sumram[28][60]+sumram[28][61]+sumram[28][62]+sumram[28][63]+sumram[28][64]+sumram[28][65]+sumram[28][66]+sumram[28][67]+sumram[28][68]+sumram[28][69]+sumram[28][70]+sumram[28][71]+sumram[28][72]+sumram[28][73]+sumram[28][74]+sumram[28][75]+sumram[28][76]+sumram[28][77]+sumram[28][78]+sumram[28][79]+sumram[28][80]+sumram[28][81]+sumram[28][82]+sumram[28][83]+sumram[28][84]+sumram[28][85]+sumram[28][86]+sumram[28][87]+sumram[28][88]+sumram[28][89]+sumram[28][90]+sumram[28][91]+sumram[28][92]+sumram[28][93]+sumram[28][94]+sumram[28][95]+sumram[28][96]+sumram[28][97]+sumram[28][98]+sumram[28][99]+sumram[28][100]+sumram[28][101]+sumram[28][102]+sumram[28][103]+sumram[28][104]+sumram[28][105]+sumram[28][106]+sumram[28][107]+sumram[28][108]+sumram[28][109]+sumram[28][110]+sumram[28][111]+sumram[28][112]+sumram[28][113]+sumram[28][114]+sumram[28][115]+sumram[28][116]+sumram[28][117]+sumram[28][118]+sumram[28][119]+sumram[28][120]+sumram[28][121]+sumram[28][122]+sumram[28][123]+sumram[28][124]+sumram[28][125]+sumram[28][126]+sumram[28][127]+sumram[28][128]+sumram[28][129]+sumram[28][130]+sumram[28][131]+sumram[28][132]+sumram[28][133]+sumram[28][134]+sumram[28][135]+sumram[28][136];
    assign sumcache[29]=sumram[29][0]+sumram[29][1]+sumram[29][2]+sumram[29][3]+sumram[29][4]+sumram[29][5]+sumram[29][6]+sumram[29][7]+sumram[29][8]+sumram[29][9]+sumram[29][10]+sumram[29][11]+sumram[29][12]+sumram[29][13]+sumram[29][14]+sumram[29][15]+sumram[29][16]+sumram[29][17]+sumram[29][18]+sumram[29][19]+sumram[29][20]+sumram[29][21]+sumram[29][22]+sumram[29][23]+sumram[29][24]+sumram[29][25]+sumram[29][26]+sumram[29][27]+sumram[29][28]+sumram[29][29]+sumram[29][30]+sumram[29][31]+sumram[29][32]+sumram[29][33]+sumram[29][34]+sumram[29][35]+sumram[29][36]+sumram[29][37]+sumram[29][38]+sumram[29][39]+sumram[29][40]+sumram[29][41]+sumram[29][42]+sumram[29][43]+sumram[29][44]+sumram[29][45]+sumram[29][46]+sumram[29][47]+sumram[29][48]+sumram[29][49]+sumram[29][50]+sumram[29][51]+sumram[29][52]+sumram[29][53]+sumram[29][54]+sumram[29][55]+sumram[29][56]+sumram[29][57]+sumram[29][58]+sumram[29][59]+sumram[29][60]+sumram[29][61]+sumram[29][62]+sumram[29][63]+sumram[29][64]+sumram[29][65]+sumram[29][66]+sumram[29][67]+sumram[29][68]+sumram[29][69]+sumram[29][70]+sumram[29][71]+sumram[29][72]+sumram[29][73]+sumram[29][74]+sumram[29][75]+sumram[29][76]+sumram[29][77]+sumram[29][78]+sumram[29][79]+sumram[29][80]+sumram[29][81]+sumram[29][82]+sumram[29][83]+sumram[29][84]+sumram[29][85]+sumram[29][86]+sumram[29][87]+sumram[29][88]+sumram[29][89]+sumram[29][90]+sumram[29][91]+sumram[29][92]+sumram[29][93]+sumram[29][94]+sumram[29][95]+sumram[29][96]+sumram[29][97]+sumram[29][98]+sumram[29][99]+sumram[29][100]+sumram[29][101]+sumram[29][102]+sumram[29][103]+sumram[29][104]+sumram[29][105]+sumram[29][106]+sumram[29][107]+sumram[29][108]+sumram[29][109]+sumram[29][110]+sumram[29][111]+sumram[29][112]+sumram[29][113]+sumram[29][114]+sumram[29][115]+sumram[29][116]+sumram[29][117]+sumram[29][118]+sumram[29][119]+sumram[29][120]+sumram[29][121]+sumram[29][122]+sumram[29][123]+sumram[29][124]+sumram[29][125]+sumram[29][126]+sumram[29][127]+sumram[29][128]+sumram[29][129]+sumram[29][130]+sumram[29][131]+sumram[29][132]+sumram[29][133]+sumram[29][134]+sumram[29][135]+sumram[29][136];
    assign sumcache[30]=sumram[30][0]+sumram[30][1]+sumram[30][2]+sumram[30][3]+sumram[30][4]+sumram[30][5]+sumram[30][6]+sumram[30][7]+sumram[30][8]+sumram[30][9]+sumram[30][10]+sumram[30][11]+sumram[30][12]+sumram[30][13]+sumram[30][14]+sumram[30][15]+sumram[30][16]+sumram[30][17]+sumram[30][18]+sumram[30][19]+sumram[30][20]+sumram[30][21]+sumram[30][22]+sumram[30][23]+sumram[30][24]+sumram[30][25]+sumram[30][26]+sumram[30][27]+sumram[30][28]+sumram[30][29]+sumram[30][30]+sumram[30][31]+sumram[30][32]+sumram[30][33]+sumram[30][34]+sumram[30][35]+sumram[30][36]+sumram[30][37]+sumram[30][38]+sumram[30][39]+sumram[30][40]+sumram[30][41]+sumram[30][42]+sumram[30][43]+sumram[30][44]+sumram[30][45]+sumram[30][46]+sumram[30][47]+sumram[30][48]+sumram[30][49]+sumram[30][50]+sumram[30][51]+sumram[30][52]+sumram[30][53]+sumram[30][54]+sumram[30][55]+sumram[30][56]+sumram[30][57]+sumram[30][58]+sumram[30][59]+sumram[30][60]+sumram[30][61]+sumram[30][62]+sumram[30][63]+sumram[30][64]+sumram[30][65]+sumram[30][66]+sumram[30][67]+sumram[30][68]+sumram[30][69]+sumram[30][70]+sumram[30][71]+sumram[30][72]+sumram[30][73]+sumram[30][74]+sumram[30][75]+sumram[30][76]+sumram[30][77]+sumram[30][78]+sumram[30][79]+sumram[30][80]+sumram[30][81]+sumram[30][82]+sumram[30][83]+sumram[30][84]+sumram[30][85]+sumram[30][86]+sumram[30][87]+sumram[30][88]+sumram[30][89]+sumram[30][90]+sumram[30][91]+sumram[30][92]+sumram[30][93]+sumram[30][94]+sumram[30][95]+sumram[30][96]+sumram[30][97]+sumram[30][98]+sumram[30][99]+sumram[30][100]+sumram[30][101]+sumram[30][102]+sumram[30][103]+sumram[30][104]+sumram[30][105]+sumram[30][106]+sumram[30][107]+sumram[30][108]+sumram[30][109]+sumram[30][110]+sumram[30][111]+sumram[30][112]+sumram[30][113]+sumram[30][114]+sumram[30][115]+sumram[30][116]+sumram[30][117]+sumram[30][118]+sumram[30][119]+sumram[30][120]+sumram[30][121]+sumram[30][122]+sumram[30][123]+sumram[30][124]+sumram[30][125]+sumram[30][126]+sumram[30][127]+sumram[30][128]+sumram[30][129]+sumram[30][130]+sumram[30][131]+sumram[30][132]+sumram[30][133]+sumram[30][134]+sumram[30][135]+sumram[30][136];
    assign sumcache[31]=sumram[31][0]+sumram[31][1]+sumram[31][2]+sumram[31][3]+sumram[31][4]+sumram[31][5]+sumram[31][6]+sumram[31][7]+sumram[31][8]+sumram[31][9]+sumram[31][10]+sumram[31][11]+sumram[31][12]+sumram[31][13]+sumram[31][14]+sumram[31][15]+sumram[31][16]+sumram[31][17]+sumram[31][18]+sumram[31][19]+sumram[31][20]+sumram[31][21]+sumram[31][22]+sumram[31][23]+sumram[31][24]+sumram[31][25]+sumram[31][26]+sumram[31][27]+sumram[31][28]+sumram[31][29]+sumram[31][30]+sumram[31][31]+sumram[31][32]+sumram[31][33]+sumram[31][34]+sumram[31][35]+sumram[31][36]+sumram[31][37]+sumram[31][38]+sumram[31][39]+sumram[31][40]+sumram[31][41]+sumram[31][42]+sumram[31][43]+sumram[31][44]+sumram[31][45]+sumram[31][46]+sumram[31][47]+sumram[31][48]+sumram[31][49]+sumram[31][50]+sumram[31][51]+sumram[31][52]+sumram[31][53]+sumram[31][54]+sumram[31][55]+sumram[31][56]+sumram[31][57]+sumram[31][58]+sumram[31][59]+sumram[31][60]+sumram[31][61]+sumram[31][62]+sumram[31][63]+sumram[31][64]+sumram[31][65]+sumram[31][66]+sumram[31][67]+sumram[31][68]+sumram[31][69]+sumram[31][70]+sumram[31][71]+sumram[31][72]+sumram[31][73]+sumram[31][74]+sumram[31][75]+sumram[31][76]+sumram[31][77]+sumram[31][78]+sumram[31][79]+sumram[31][80]+sumram[31][81]+sumram[31][82]+sumram[31][83]+sumram[31][84]+sumram[31][85]+sumram[31][86]+sumram[31][87]+sumram[31][88]+sumram[31][89]+sumram[31][90]+sumram[31][91]+sumram[31][92]+sumram[31][93]+sumram[31][94]+sumram[31][95]+sumram[31][96]+sumram[31][97]+sumram[31][98]+sumram[31][99]+sumram[31][100]+sumram[31][101]+sumram[31][102]+sumram[31][103]+sumram[31][104]+sumram[31][105]+sumram[31][106]+sumram[31][107]+sumram[31][108]+sumram[31][109]+sumram[31][110]+sumram[31][111]+sumram[31][112]+sumram[31][113]+sumram[31][114]+sumram[31][115]+sumram[31][116]+sumram[31][117]+sumram[31][118]+sumram[31][119]+sumram[31][120]+sumram[31][121]+sumram[31][122]+sumram[31][123]+sumram[31][124]+sumram[31][125]+sumram[31][126]+sumram[31][127]+sumram[31][128]+sumram[31][129]+sumram[31][130]+sumram[31][131]+sumram[31][132]+sumram[31][133]+sumram[31][134]+sumram[31][135]+sumram[31][136];
    assign sumcache[32]=sumram[32][0]+sumram[32][1]+sumram[32][2]+sumram[32][3]+sumram[32][4]+sumram[32][5]+sumram[32][6]+sumram[32][7]+sumram[32][8]+sumram[32][9]+sumram[32][10]+sumram[32][11]+sumram[32][12]+sumram[32][13]+sumram[32][14]+sumram[32][15]+sumram[32][16]+sumram[32][17]+sumram[32][18]+sumram[32][19]+sumram[32][20]+sumram[32][21]+sumram[32][22]+sumram[32][23]+sumram[32][24]+sumram[32][25]+sumram[32][26]+sumram[32][27]+sumram[32][28]+sumram[32][29]+sumram[32][30]+sumram[32][31]+sumram[32][32]+sumram[32][33]+sumram[32][34]+sumram[32][35]+sumram[32][36]+sumram[32][37]+sumram[32][38]+sumram[32][39]+sumram[32][40]+sumram[32][41]+sumram[32][42]+sumram[32][43]+sumram[32][44]+sumram[32][45]+sumram[32][46]+sumram[32][47]+sumram[32][48]+sumram[32][49]+sumram[32][50]+sumram[32][51]+sumram[32][52]+sumram[32][53]+sumram[32][54]+sumram[32][55]+sumram[32][56]+sumram[32][57]+sumram[32][58]+sumram[32][59]+sumram[32][60]+sumram[32][61]+sumram[32][62]+sumram[32][63]+sumram[32][64]+sumram[32][65]+sumram[32][66]+sumram[32][67]+sumram[32][68]+sumram[32][69]+sumram[32][70]+sumram[32][71]+sumram[32][72]+sumram[32][73]+sumram[32][74]+sumram[32][75]+sumram[32][76]+sumram[32][77]+sumram[32][78]+sumram[32][79]+sumram[32][80]+sumram[32][81]+sumram[32][82]+sumram[32][83]+sumram[32][84]+sumram[32][85]+sumram[32][86]+sumram[32][87]+sumram[32][88]+sumram[32][89]+sumram[32][90]+sumram[32][91]+sumram[32][92]+sumram[32][93]+sumram[32][94]+sumram[32][95]+sumram[32][96]+sumram[32][97]+sumram[32][98]+sumram[32][99]+sumram[32][100]+sumram[32][101]+sumram[32][102]+sumram[32][103]+sumram[32][104]+sumram[32][105]+sumram[32][106]+sumram[32][107]+sumram[32][108]+sumram[32][109]+sumram[32][110]+sumram[32][111]+sumram[32][112]+sumram[32][113]+sumram[32][114]+sumram[32][115]+sumram[32][116]+sumram[32][117]+sumram[32][118]+sumram[32][119]+sumram[32][120]+sumram[32][121]+sumram[32][122]+sumram[32][123]+sumram[32][124]+sumram[32][125]+sumram[32][126]+sumram[32][127]+sumram[32][128]+sumram[32][129]+sumram[32][130]+sumram[32][131]+sumram[32][132]+sumram[32][133]+sumram[32][134]+sumram[32][135]+sumram[32][136];
    assign sumcache[33]=sumram[33][0]+sumram[33][1]+sumram[33][2]+sumram[33][3]+sumram[33][4]+sumram[33][5]+sumram[33][6]+sumram[33][7]+sumram[33][8]+sumram[33][9]+sumram[33][10]+sumram[33][11]+sumram[33][12]+sumram[33][13]+sumram[33][14]+sumram[33][15]+sumram[33][16]+sumram[33][17]+sumram[33][18]+sumram[33][19]+sumram[33][20]+sumram[33][21]+sumram[33][22]+sumram[33][23]+sumram[33][24]+sumram[33][25]+sumram[33][26]+sumram[33][27]+sumram[33][28]+sumram[33][29]+sumram[33][30]+sumram[33][31]+sumram[33][32]+sumram[33][33]+sumram[33][34]+sumram[33][35]+sumram[33][36]+sumram[33][37]+sumram[33][38]+sumram[33][39]+sumram[33][40]+sumram[33][41]+sumram[33][42]+sumram[33][43]+sumram[33][44]+sumram[33][45]+sumram[33][46]+sumram[33][47]+sumram[33][48]+sumram[33][49]+sumram[33][50]+sumram[33][51]+sumram[33][52]+sumram[33][53]+sumram[33][54]+sumram[33][55]+sumram[33][56]+sumram[33][57]+sumram[33][58]+sumram[33][59]+sumram[33][60]+sumram[33][61]+sumram[33][62]+sumram[33][63]+sumram[33][64]+sumram[33][65]+sumram[33][66]+sumram[33][67]+sumram[33][68]+sumram[33][69]+sumram[33][70]+sumram[33][71]+sumram[33][72]+sumram[33][73]+sumram[33][74]+sumram[33][75]+sumram[33][76]+sumram[33][77]+sumram[33][78]+sumram[33][79]+sumram[33][80]+sumram[33][81]+sumram[33][82]+sumram[33][83]+sumram[33][84]+sumram[33][85]+sumram[33][86]+sumram[33][87]+sumram[33][88]+sumram[33][89]+sumram[33][90]+sumram[33][91]+sumram[33][92]+sumram[33][93]+sumram[33][94]+sumram[33][95]+sumram[33][96]+sumram[33][97]+sumram[33][98]+sumram[33][99]+sumram[33][100]+sumram[33][101]+sumram[33][102]+sumram[33][103]+sumram[33][104]+sumram[33][105]+sumram[33][106]+sumram[33][107]+sumram[33][108]+sumram[33][109]+sumram[33][110]+sumram[33][111]+sumram[33][112]+sumram[33][113]+sumram[33][114]+sumram[33][115]+sumram[33][116]+sumram[33][117]+sumram[33][118]+sumram[33][119]+sumram[33][120]+sumram[33][121]+sumram[33][122]+sumram[33][123]+sumram[33][124]+sumram[33][125]+sumram[33][126]+sumram[33][127]+sumram[33][128]+sumram[33][129]+sumram[33][130]+sumram[33][131]+sumram[33][132]+sumram[33][133]+sumram[33][134]+sumram[33][135]+sumram[33][136];
    assign sumcache[34]=sumram[34][0]+sumram[34][1]+sumram[34][2]+sumram[34][3]+sumram[34][4]+sumram[34][5]+sumram[34][6]+sumram[34][7]+sumram[34][8]+sumram[34][9]+sumram[34][10]+sumram[34][11]+sumram[34][12]+sumram[34][13]+sumram[34][14]+sumram[34][15]+sumram[34][16]+sumram[34][17]+sumram[34][18]+sumram[34][19]+sumram[34][20]+sumram[34][21]+sumram[34][22]+sumram[34][23]+sumram[34][24]+sumram[34][25]+sumram[34][26]+sumram[34][27]+sumram[34][28]+sumram[34][29]+sumram[34][30]+sumram[34][31]+sumram[34][32]+sumram[34][33]+sumram[34][34]+sumram[34][35]+sumram[34][36]+sumram[34][37]+sumram[34][38]+sumram[34][39]+sumram[34][40]+sumram[34][41]+sumram[34][42]+sumram[34][43]+sumram[34][44]+sumram[34][45]+sumram[34][46]+sumram[34][47]+sumram[34][48]+sumram[34][49]+sumram[34][50]+sumram[34][51]+sumram[34][52]+sumram[34][53]+sumram[34][54]+sumram[34][55]+sumram[34][56]+sumram[34][57]+sumram[34][58]+sumram[34][59]+sumram[34][60]+sumram[34][61]+sumram[34][62]+sumram[34][63]+sumram[34][64]+sumram[34][65]+sumram[34][66]+sumram[34][67]+sumram[34][68]+sumram[34][69]+sumram[34][70]+sumram[34][71]+sumram[34][72]+sumram[34][73]+sumram[34][74]+sumram[34][75]+sumram[34][76]+sumram[34][77]+sumram[34][78]+sumram[34][79]+sumram[34][80]+sumram[34][81]+sumram[34][82]+sumram[34][83]+sumram[34][84]+sumram[34][85]+sumram[34][86]+sumram[34][87]+sumram[34][88]+sumram[34][89]+sumram[34][90]+sumram[34][91]+sumram[34][92]+sumram[34][93]+sumram[34][94]+sumram[34][95]+sumram[34][96]+sumram[34][97]+sumram[34][98]+sumram[34][99]+sumram[34][100]+sumram[34][101]+sumram[34][102]+sumram[34][103]+sumram[34][104]+sumram[34][105]+sumram[34][106]+sumram[34][107]+sumram[34][108]+sumram[34][109]+sumram[34][110]+sumram[34][111]+sumram[34][112]+sumram[34][113]+sumram[34][114]+sumram[34][115]+sumram[34][116]+sumram[34][117]+sumram[34][118]+sumram[34][119]+sumram[34][120]+sumram[34][121]+sumram[34][122]+sumram[34][123]+sumram[34][124]+sumram[34][125]+sumram[34][126]+sumram[34][127]+sumram[34][128]+sumram[34][129]+sumram[34][130]+sumram[34][131]+sumram[34][132]+sumram[34][133]+sumram[34][134]+sumram[34][135]+sumram[34][136];
    assign sumcache[35]=sumram[35][0]+sumram[35][1]+sumram[35][2]+sumram[35][3]+sumram[35][4]+sumram[35][5]+sumram[35][6]+sumram[35][7]+sumram[35][8]+sumram[35][9]+sumram[35][10]+sumram[35][11]+sumram[35][12]+sumram[35][13]+sumram[35][14]+sumram[35][15]+sumram[35][16]+sumram[35][17]+sumram[35][18]+sumram[35][19]+sumram[35][20]+sumram[35][21]+sumram[35][22]+sumram[35][23]+sumram[35][24]+sumram[35][25]+sumram[35][26]+sumram[35][27]+sumram[35][28]+sumram[35][29]+sumram[35][30]+sumram[35][31]+sumram[35][32]+sumram[35][33]+sumram[35][34]+sumram[35][35]+sumram[35][36]+sumram[35][37]+sumram[35][38]+sumram[35][39]+sumram[35][40]+sumram[35][41]+sumram[35][42]+sumram[35][43]+sumram[35][44]+sumram[35][45]+sumram[35][46]+sumram[35][47]+sumram[35][48]+sumram[35][49]+sumram[35][50]+sumram[35][51]+sumram[35][52]+sumram[35][53]+sumram[35][54]+sumram[35][55]+sumram[35][56]+sumram[35][57]+sumram[35][58]+sumram[35][59]+sumram[35][60]+sumram[35][61]+sumram[35][62]+sumram[35][63]+sumram[35][64]+sumram[35][65]+sumram[35][66]+sumram[35][67]+sumram[35][68]+sumram[35][69]+sumram[35][70]+sumram[35][71]+sumram[35][72]+sumram[35][73]+sumram[35][74]+sumram[35][75]+sumram[35][76]+sumram[35][77]+sumram[35][78]+sumram[35][79]+sumram[35][80]+sumram[35][81]+sumram[35][82]+sumram[35][83]+sumram[35][84]+sumram[35][85]+sumram[35][86]+sumram[35][87]+sumram[35][88]+sumram[35][89]+sumram[35][90]+sumram[35][91]+sumram[35][92]+sumram[35][93]+sumram[35][94]+sumram[35][95]+sumram[35][96]+sumram[35][97]+sumram[35][98]+sumram[35][99]+sumram[35][100]+sumram[35][101]+sumram[35][102]+sumram[35][103]+sumram[35][104]+sumram[35][105]+sumram[35][106]+sumram[35][107]+sumram[35][108]+sumram[35][109]+sumram[35][110]+sumram[35][111]+sumram[35][112]+sumram[35][113]+sumram[35][114]+sumram[35][115]+sumram[35][116]+sumram[35][117]+sumram[35][118]+sumram[35][119]+sumram[35][120]+sumram[35][121]+sumram[35][122]+sumram[35][123]+sumram[35][124]+sumram[35][125]+sumram[35][126]+sumram[35][127]+sumram[35][128]+sumram[35][129]+sumram[35][130]+sumram[35][131]+sumram[35][132]+sumram[35][133]+sumram[35][134]+sumram[35][135]+sumram[35][136];
    assign sumcache[36]=sumram[36][0]+sumram[36][1]+sumram[36][2]+sumram[36][3]+sumram[36][4]+sumram[36][5]+sumram[36][6]+sumram[36][7]+sumram[36][8]+sumram[36][9]+sumram[36][10]+sumram[36][11]+sumram[36][12]+sumram[36][13]+sumram[36][14]+sumram[36][15]+sumram[36][16]+sumram[36][17]+sumram[36][18]+sumram[36][19]+sumram[36][20]+sumram[36][21]+sumram[36][22]+sumram[36][23]+sumram[36][24]+sumram[36][25]+sumram[36][26]+sumram[36][27]+sumram[36][28]+sumram[36][29]+sumram[36][30]+sumram[36][31]+sumram[36][32]+sumram[36][33]+sumram[36][34]+sumram[36][35]+sumram[36][36]+sumram[36][37]+sumram[36][38]+sumram[36][39]+sumram[36][40]+sumram[36][41]+sumram[36][42]+sumram[36][43]+sumram[36][44]+sumram[36][45]+sumram[36][46]+sumram[36][47]+sumram[36][48]+sumram[36][49]+sumram[36][50]+sumram[36][51]+sumram[36][52]+sumram[36][53]+sumram[36][54]+sumram[36][55]+sumram[36][56]+sumram[36][57]+sumram[36][58]+sumram[36][59]+sumram[36][60]+sumram[36][61]+sumram[36][62]+sumram[36][63]+sumram[36][64]+sumram[36][65]+sumram[36][66]+sumram[36][67]+sumram[36][68]+sumram[36][69]+sumram[36][70]+sumram[36][71]+sumram[36][72]+sumram[36][73]+sumram[36][74]+sumram[36][75]+sumram[36][76]+sumram[36][77]+sumram[36][78]+sumram[36][79]+sumram[36][80]+sumram[36][81]+sumram[36][82]+sumram[36][83]+sumram[36][84]+sumram[36][85]+sumram[36][86]+sumram[36][87]+sumram[36][88]+sumram[36][89]+sumram[36][90]+sumram[36][91]+sumram[36][92]+sumram[36][93]+sumram[36][94]+sumram[36][95]+sumram[36][96]+sumram[36][97]+sumram[36][98]+sumram[36][99]+sumram[36][100]+sumram[36][101]+sumram[36][102]+sumram[36][103]+sumram[36][104]+sumram[36][105]+sumram[36][106]+sumram[36][107]+sumram[36][108]+sumram[36][109]+sumram[36][110]+sumram[36][111]+sumram[36][112]+sumram[36][113]+sumram[36][114]+sumram[36][115]+sumram[36][116]+sumram[36][117]+sumram[36][118]+sumram[36][119]+sumram[36][120]+sumram[36][121]+sumram[36][122]+sumram[36][123]+sumram[36][124]+sumram[36][125]+sumram[36][126]+sumram[36][127]+sumram[36][128]+sumram[36][129]+sumram[36][130]+sumram[36][131]+sumram[36][132]+sumram[36][133]+sumram[36][134]+sumram[36][135]+sumram[36][136];
    assign sumcache[37]=sumram[37][0]+sumram[37][1]+sumram[37][2]+sumram[37][3]+sumram[37][4]+sumram[37][5]+sumram[37][6]+sumram[37][7]+sumram[37][8]+sumram[37][9]+sumram[37][10]+sumram[37][11]+sumram[37][12]+sumram[37][13]+sumram[37][14]+sumram[37][15]+sumram[37][16]+sumram[37][17]+sumram[37][18]+sumram[37][19]+sumram[37][20]+sumram[37][21]+sumram[37][22]+sumram[37][23]+sumram[37][24]+sumram[37][25]+sumram[37][26]+sumram[37][27]+sumram[37][28]+sumram[37][29]+sumram[37][30]+sumram[37][31]+sumram[37][32]+sumram[37][33]+sumram[37][34]+sumram[37][35]+sumram[37][36]+sumram[37][37]+sumram[37][38]+sumram[37][39]+sumram[37][40]+sumram[37][41]+sumram[37][42]+sumram[37][43]+sumram[37][44]+sumram[37][45]+sumram[37][46]+sumram[37][47]+sumram[37][48]+sumram[37][49]+sumram[37][50]+sumram[37][51]+sumram[37][52]+sumram[37][53]+sumram[37][54]+sumram[37][55]+sumram[37][56]+sumram[37][57]+sumram[37][58]+sumram[37][59]+sumram[37][60]+sumram[37][61]+sumram[37][62]+sumram[37][63]+sumram[37][64]+sumram[37][65]+sumram[37][66]+sumram[37][67]+sumram[37][68]+sumram[37][69]+sumram[37][70]+sumram[37][71]+sumram[37][72]+sumram[37][73]+sumram[37][74]+sumram[37][75]+sumram[37][76]+sumram[37][77]+sumram[37][78]+sumram[37][79]+sumram[37][80]+sumram[37][81]+sumram[37][82]+sumram[37][83]+sumram[37][84]+sumram[37][85]+sumram[37][86]+sumram[37][87]+sumram[37][88]+sumram[37][89]+sumram[37][90]+sumram[37][91]+sumram[37][92]+sumram[37][93]+sumram[37][94]+sumram[37][95]+sumram[37][96]+sumram[37][97]+sumram[37][98]+sumram[37][99]+sumram[37][100]+sumram[37][101]+sumram[37][102]+sumram[37][103]+sumram[37][104]+sumram[37][105]+sumram[37][106]+sumram[37][107]+sumram[37][108]+sumram[37][109]+sumram[37][110]+sumram[37][111]+sumram[37][112]+sumram[37][113]+sumram[37][114]+sumram[37][115]+sumram[37][116]+sumram[37][117]+sumram[37][118]+sumram[37][119]+sumram[37][120]+sumram[37][121]+sumram[37][122]+sumram[37][123]+sumram[37][124]+sumram[37][125]+sumram[37][126]+sumram[37][127]+sumram[37][128]+sumram[37][129]+sumram[37][130]+sumram[37][131]+sumram[37][132]+sumram[37][133]+sumram[37][134]+sumram[37][135]+sumram[37][136];
    assign sumcache[38]=sumram[38][0]+sumram[38][1]+sumram[38][2]+sumram[38][3]+sumram[38][4]+sumram[38][5]+sumram[38][6]+sumram[38][7]+sumram[38][8]+sumram[38][9]+sumram[38][10]+sumram[38][11]+sumram[38][12]+sumram[38][13]+sumram[38][14]+sumram[38][15]+sumram[38][16]+sumram[38][17]+sumram[38][18]+sumram[38][19]+sumram[38][20]+sumram[38][21]+sumram[38][22]+sumram[38][23]+sumram[38][24]+sumram[38][25]+sumram[38][26]+sumram[38][27]+sumram[38][28]+sumram[38][29]+sumram[38][30]+sumram[38][31]+sumram[38][32]+sumram[38][33]+sumram[38][34]+sumram[38][35]+sumram[38][36]+sumram[38][37]+sumram[38][38]+sumram[38][39]+sumram[38][40]+sumram[38][41]+sumram[38][42]+sumram[38][43]+sumram[38][44]+sumram[38][45]+sumram[38][46]+sumram[38][47]+sumram[38][48]+sumram[38][49]+sumram[38][50]+sumram[38][51]+sumram[38][52]+sumram[38][53]+sumram[38][54]+sumram[38][55]+sumram[38][56]+sumram[38][57]+sumram[38][58]+sumram[38][59]+sumram[38][60]+sumram[38][61]+sumram[38][62]+sumram[38][63]+sumram[38][64]+sumram[38][65]+sumram[38][66]+sumram[38][67]+sumram[38][68]+sumram[38][69]+sumram[38][70]+sumram[38][71]+sumram[38][72]+sumram[38][73]+sumram[38][74]+sumram[38][75]+sumram[38][76]+sumram[38][77]+sumram[38][78]+sumram[38][79]+sumram[38][80]+sumram[38][81]+sumram[38][82]+sumram[38][83]+sumram[38][84]+sumram[38][85]+sumram[38][86]+sumram[38][87]+sumram[38][88]+sumram[38][89]+sumram[38][90]+sumram[38][91]+sumram[38][92]+sumram[38][93]+sumram[38][94]+sumram[38][95]+sumram[38][96]+sumram[38][97]+sumram[38][98]+sumram[38][99]+sumram[38][100]+sumram[38][101]+sumram[38][102]+sumram[38][103]+sumram[38][104]+sumram[38][105]+sumram[38][106]+sumram[38][107]+sumram[38][108]+sumram[38][109]+sumram[38][110]+sumram[38][111]+sumram[38][112]+sumram[38][113]+sumram[38][114]+sumram[38][115]+sumram[38][116]+sumram[38][117]+sumram[38][118]+sumram[38][119]+sumram[38][120]+sumram[38][121]+sumram[38][122]+sumram[38][123]+sumram[38][124]+sumram[38][125]+sumram[38][126]+sumram[38][127]+sumram[38][128]+sumram[38][129]+sumram[38][130]+sumram[38][131]+sumram[38][132]+sumram[38][133]+sumram[38][134]+sumram[38][135]+sumram[38][136];
    assign sumcache[39]=sumram[39][0]+sumram[39][1]+sumram[39][2]+sumram[39][3]+sumram[39][4]+sumram[39][5]+sumram[39][6]+sumram[39][7]+sumram[39][8]+sumram[39][9]+sumram[39][10]+sumram[39][11]+sumram[39][12]+sumram[39][13]+sumram[39][14]+sumram[39][15]+sumram[39][16]+sumram[39][17]+sumram[39][18]+sumram[39][19]+sumram[39][20]+sumram[39][21]+sumram[39][22]+sumram[39][23]+sumram[39][24]+sumram[39][25]+sumram[39][26]+sumram[39][27]+sumram[39][28]+sumram[39][29]+sumram[39][30]+sumram[39][31]+sumram[39][32]+sumram[39][33]+sumram[39][34]+sumram[39][35]+sumram[39][36]+sumram[39][37]+sumram[39][38]+sumram[39][39]+sumram[39][40]+sumram[39][41]+sumram[39][42]+sumram[39][43]+sumram[39][44]+sumram[39][45]+sumram[39][46]+sumram[39][47]+sumram[39][48]+sumram[39][49]+sumram[39][50]+sumram[39][51]+sumram[39][52]+sumram[39][53]+sumram[39][54]+sumram[39][55]+sumram[39][56]+sumram[39][57]+sumram[39][58]+sumram[39][59]+sumram[39][60]+sumram[39][61]+sumram[39][62]+sumram[39][63]+sumram[39][64]+sumram[39][65]+sumram[39][66]+sumram[39][67]+sumram[39][68]+sumram[39][69]+sumram[39][70]+sumram[39][71]+sumram[39][72]+sumram[39][73]+sumram[39][74]+sumram[39][75]+sumram[39][76]+sumram[39][77]+sumram[39][78]+sumram[39][79]+sumram[39][80]+sumram[39][81]+sumram[39][82]+sumram[39][83]+sumram[39][84]+sumram[39][85]+sumram[39][86]+sumram[39][87]+sumram[39][88]+sumram[39][89]+sumram[39][90]+sumram[39][91]+sumram[39][92]+sumram[39][93]+sumram[39][94]+sumram[39][95]+sumram[39][96]+sumram[39][97]+sumram[39][98]+sumram[39][99]+sumram[39][100]+sumram[39][101]+sumram[39][102]+sumram[39][103]+sumram[39][104]+sumram[39][105]+sumram[39][106]+sumram[39][107]+sumram[39][108]+sumram[39][109]+sumram[39][110]+sumram[39][111]+sumram[39][112]+sumram[39][113]+sumram[39][114]+sumram[39][115]+sumram[39][116]+sumram[39][117]+sumram[39][118]+sumram[39][119]+sumram[39][120]+sumram[39][121]+sumram[39][122]+sumram[39][123]+sumram[39][124]+sumram[39][125]+sumram[39][126]+sumram[39][127]+sumram[39][128]+sumram[39][129]+sumram[39][130]+sumram[39][131]+sumram[39][132]+sumram[39][133]+sumram[39][134]+sumram[39][135]+sumram[39][136];
    assign sumcache[40]=sumram[40][0]+sumram[40][1]+sumram[40][2]+sumram[40][3]+sumram[40][4]+sumram[40][5]+sumram[40][6]+sumram[40][7]+sumram[40][8]+sumram[40][9]+sumram[40][10]+sumram[40][11]+sumram[40][12]+sumram[40][13]+sumram[40][14]+sumram[40][15]+sumram[40][16]+sumram[40][17]+sumram[40][18]+sumram[40][19]+sumram[40][20]+sumram[40][21]+sumram[40][22]+sumram[40][23]+sumram[40][24]+sumram[40][25]+sumram[40][26]+sumram[40][27]+sumram[40][28]+sumram[40][29]+sumram[40][30]+sumram[40][31]+sumram[40][32]+sumram[40][33]+sumram[40][34]+sumram[40][35]+sumram[40][36]+sumram[40][37]+sumram[40][38]+sumram[40][39]+sumram[40][40]+sumram[40][41]+sumram[40][42]+sumram[40][43]+sumram[40][44]+sumram[40][45]+sumram[40][46]+sumram[40][47]+sumram[40][48]+sumram[40][49]+sumram[40][50]+sumram[40][51]+sumram[40][52]+sumram[40][53]+sumram[40][54]+sumram[40][55]+sumram[40][56]+sumram[40][57]+sumram[40][58]+sumram[40][59]+sumram[40][60]+sumram[40][61]+sumram[40][62]+sumram[40][63]+sumram[40][64]+sumram[40][65]+sumram[40][66]+sumram[40][67]+sumram[40][68]+sumram[40][69]+sumram[40][70]+sumram[40][71]+sumram[40][72]+sumram[40][73]+sumram[40][74]+sumram[40][75]+sumram[40][76]+sumram[40][77]+sumram[40][78]+sumram[40][79]+sumram[40][80]+sumram[40][81]+sumram[40][82]+sumram[40][83]+sumram[40][84]+sumram[40][85]+sumram[40][86]+sumram[40][87]+sumram[40][88]+sumram[40][89]+sumram[40][90]+sumram[40][91]+sumram[40][92]+sumram[40][93]+sumram[40][94]+sumram[40][95]+sumram[40][96]+sumram[40][97]+sumram[40][98]+sumram[40][99]+sumram[40][100]+sumram[40][101]+sumram[40][102]+sumram[40][103]+sumram[40][104]+sumram[40][105]+sumram[40][106]+sumram[40][107]+sumram[40][108]+sumram[40][109]+sumram[40][110]+sumram[40][111]+sumram[40][112]+sumram[40][113]+sumram[40][114]+sumram[40][115]+sumram[40][116]+sumram[40][117]+sumram[40][118]+sumram[40][119]+sumram[40][120]+sumram[40][121]+sumram[40][122]+sumram[40][123]+sumram[40][124]+sumram[40][125]+sumram[40][126]+sumram[40][127]+sumram[40][128]+sumram[40][129]+sumram[40][130]+sumram[40][131]+sumram[40][132]+sumram[40][133]+sumram[40][134]+sumram[40][135]+sumram[40][136];
    assign sumcache[41]=sumram[41][0]+sumram[41][1]+sumram[41][2]+sumram[41][3]+sumram[41][4]+sumram[41][5]+sumram[41][6]+sumram[41][7]+sumram[41][8]+sumram[41][9]+sumram[41][10]+sumram[41][11]+sumram[41][12]+sumram[41][13]+sumram[41][14]+sumram[41][15]+sumram[41][16]+sumram[41][17]+sumram[41][18]+sumram[41][19]+sumram[41][20]+sumram[41][21]+sumram[41][22]+sumram[41][23]+sumram[41][24]+sumram[41][25]+sumram[41][26]+sumram[41][27]+sumram[41][28]+sumram[41][29]+sumram[41][30]+sumram[41][31]+sumram[41][32]+sumram[41][33]+sumram[41][34]+sumram[41][35]+sumram[41][36]+sumram[41][37]+sumram[41][38]+sumram[41][39]+sumram[41][40]+sumram[41][41]+sumram[41][42]+sumram[41][43]+sumram[41][44]+sumram[41][45]+sumram[41][46]+sumram[41][47]+sumram[41][48]+sumram[41][49]+sumram[41][50]+sumram[41][51]+sumram[41][52]+sumram[41][53]+sumram[41][54]+sumram[41][55]+sumram[41][56]+sumram[41][57]+sumram[41][58]+sumram[41][59]+sumram[41][60]+sumram[41][61]+sumram[41][62]+sumram[41][63]+sumram[41][64]+sumram[41][65]+sumram[41][66]+sumram[41][67]+sumram[41][68]+sumram[41][69]+sumram[41][70]+sumram[41][71]+sumram[41][72]+sumram[41][73]+sumram[41][74]+sumram[41][75]+sumram[41][76]+sumram[41][77]+sumram[41][78]+sumram[41][79]+sumram[41][80]+sumram[41][81]+sumram[41][82]+sumram[41][83]+sumram[41][84]+sumram[41][85]+sumram[41][86]+sumram[41][87]+sumram[41][88]+sumram[41][89]+sumram[41][90]+sumram[41][91]+sumram[41][92]+sumram[41][93]+sumram[41][94]+sumram[41][95]+sumram[41][96]+sumram[41][97]+sumram[41][98]+sumram[41][99]+sumram[41][100]+sumram[41][101]+sumram[41][102]+sumram[41][103]+sumram[41][104]+sumram[41][105]+sumram[41][106]+sumram[41][107]+sumram[41][108]+sumram[41][109]+sumram[41][110]+sumram[41][111]+sumram[41][112]+sumram[41][113]+sumram[41][114]+sumram[41][115]+sumram[41][116]+sumram[41][117]+sumram[41][118]+sumram[41][119]+sumram[41][120]+sumram[41][121]+sumram[41][122]+sumram[41][123]+sumram[41][124]+sumram[41][125]+sumram[41][126]+sumram[41][127]+sumram[41][128]+sumram[41][129]+sumram[41][130]+sumram[41][131]+sumram[41][132]+sumram[41][133]+sumram[41][134]+sumram[41][135]+sumram[41][136];
    assign sumcache[42]=sumram[42][0]+sumram[42][1]+sumram[42][2]+sumram[42][3]+sumram[42][4]+sumram[42][5]+sumram[42][6]+sumram[42][7]+sumram[42][8]+sumram[42][9]+sumram[42][10]+sumram[42][11]+sumram[42][12]+sumram[42][13]+sumram[42][14]+sumram[42][15]+sumram[42][16]+sumram[42][17]+sumram[42][18]+sumram[42][19]+sumram[42][20]+sumram[42][21]+sumram[42][22]+sumram[42][23]+sumram[42][24]+sumram[42][25]+sumram[42][26]+sumram[42][27]+sumram[42][28]+sumram[42][29]+sumram[42][30]+sumram[42][31]+sumram[42][32]+sumram[42][33]+sumram[42][34]+sumram[42][35]+sumram[42][36]+sumram[42][37]+sumram[42][38]+sumram[42][39]+sumram[42][40]+sumram[42][41]+sumram[42][42]+sumram[42][43]+sumram[42][44]+sumram[42][45]+sumram[42][46]+sumram[42][47]+sumram[42][48]+sumram[42][49]+sumram[42][50]+sumram[42][51]+sumram[42][52]+sumram[42][53]+sumram[42][54]+sumram[42][55]+sumram[42][56]+sumram[42][57]+sumram[42][58]+sumram[42][59]+sumram[42][60]+sumram[42][61]+sumram[42][62]+sumram[42][63]+sumram[42][64]+sumram[42][65]+sumram[42][66]+sumram[42][67]+sumram[42][68]+sumram[42][69]+sumram[42][70]+sumram[42][71]+sumram[42][72]+sumram[42][73]+sumram[42][74]+sumram[42][75]+sumram[42][76]+sumram[42][77]+sumram[42][78]+sumram[42][79]+sumram[42][80]+sumram[42][81]+sumram[42][82]+sumram[42][83]+sumram[42][84]+sumram[42][85]+sumram[42][86]+sumram[42][87]+sumram[42][88]+sumram[42][89]+sumram[42][90]+sumram[42][91]+sumram[42][92]+sumram[42][93]+sumram[42][94]+sumram[42][95]+sumram[42][96]+sumram[42][97]+sumram[42][98]+sumram[42][99]+sumram[42][100]+sumram[42][101]+sumram[42][102]+sumram[42][103]+sumram[42][104]+sumram[42][105]+sumram[42][106]+sumram[42][107]+sumram[42][108]+sumram[42][109]+sumram[42][110]+sumram[42][111]+sumram[42][112]+sumram[42][113]+sumram[42][114]+sumram[42][115]+sumram[42][116]+sumram[42][117]+sumram[42][118]+sumram[42][119]+sumram[42][120]+sumram[42][121]+sumram[42][122]+sumram[42][123]+sumram[42][124]+sumram[42][125]+sumram[42][126]+sumram[42][127]+sumram[42][128]+sumram[42][129]+sumram[42][130]+sumram[42][131]+sumram[42][132]+sumram[42][133]+sumram[42][134]+sumram[42][135]+sumram[42][136];
    assign sumcache[43]=sumram[43][0]+sumram[43][1]+sumram[43][2]+sumram[43][3]+sumram[43][4]+sumram[43][5]+sumram[43][6]+sumram[43][7]+sumram[43][8]+sumram[43][9]+sumram[43][10]+sumram[43][11]+sumram[43][12]+sumram[43][13]+sumram[43][14]+sumram[43][15]+sumram[43][16]+sumram[43][17]+sumram[43][18]+sumram[43][19]+sumram[43][20]+sumram[43][21]+sumram[43][22]+sumram[43][23]+sumram[43][24]+sumram[43][25]+sumram[43][26]+sumram[43][27]+sumram[43][28]+sumram[43][29]+sumram[43][30]+sumram[43][31]+sumram[43][32]+sumram[43][33]+sumram[43][34]+sumram[43][35]+sumram[43][36]+sumram[43][37]+sumram[43][38]+sumram[43][39]+sumram[43][40]+sumram[43][41]+sumram[43][42]+sumram[43][43]+sumram[43][44]+sumram[43][45]+sumram[43][46]+sumram[43][47]+sumram[43][48]+sumram[43][49]+sumram[43][50]+sumram[43][51]+sumram[43][52]+sumram[43][53]+sumram[43][54]+sumram[43][55]+sumram[43][56]+sumram[43][57]+sumram[43][58]+sumram[43][59]+sumram[43][60]+sumram[43][61]+sumram[43][62]+sumram[43][63]+sumram[43][64]+sumram[43][65]+sumram[43][66]+sumram[43][67]+sumram[43][68]+sumram[43][69]+sumram[43][70]+sumram[43][71]+sumram[43][72]+sumram[43][73]+sumram[43][74]+sumram[43][75]+sumram[43][76]+sumram[43][77]+sumram[43][78]+sumram[43][79]+sumram[43][80]+sumram[43][81]+sumram[43][82]+sumram[43][83]+sumram[43][84]+sumram[43][85]+sumram[43][86]+sumram[43][87]+sumram[43][88]+sumram[43][89]+sumram[43][90]+sumram[43][91]+sumram[43][92]+sumram[43][93]+sumram[43][94]+sumram[43][95]+sumram[43][96]+sumram[43][97]+sumram[43][98]+sumram[43][99]+sumram[43][100]+sumram[43][101]+sumram[43][102]+sumram[43][103]+sumram[43][104]+sumram[43][105]+sumram[43][106]+sumram[43][107]+sumram[43][108]+sumram[43][109]+sumram[43][110]+sumram[43][111]+sumram[43][112]+sumram[43][113]+sumram[43][114]+sumram[43][115]+sumram[43][116]+sumram[43][117]+sumram[43][118]+sumram[43][119]+sumram[43][120]+sumram[43][121]+sumram[43][122]+sumram[43][123]+sumram[43][124]+sumram[43][125]+sumram[43][126]+sumram[43][127]+sumram[43][128]+sumram[43][129]+sumram[43][130]+sumram[43][131]+sumram[43][132]+sumram[43][133]+sumram[43][134]+sumram[43][135]+sumram[43][136];
    assign sumcache[44]=sumram[44][0]+sumram[44][1]+sumram[44][2]+sumram[44][3]+sumram[44][4]+sumram[44][5]+sumram[44][6]+sumram[44][7]+sumram[44][8]+sumram[44][9]+sumram[44][10]+sumram[44][11]+sumram[44][12]+sumram[44][13]+sumram[44][14]+sumram[44][15]+sumram[44][16]+sumram[44][17]+sumram[44][18]+sumram[44][19]+sumram[44][20]+sumram[44][21]+sumram[44][22]+sumram[44][23]+sumram[44][24]+sumram[44][25]+sumram[44][26]+sumram[44][27]+sumram[44][28]+sumram[44][29]+sumram[44][30]+sumram[44][31]+sumram[44][32]+sumram[44][33]+sumram[44][34]+sumram[44][35]+sumram[44][36]+sumram[44][37]+sumram[44][38]+sumram[44][39]+sumram[44][40]+sumram[44][41]+sumram[44][42]+sumram[44][43]+sumram[44][44]+sumram[44][45]+sumram[44][46]+sumram[44][47]+sumram[44][48]+sumram[44][49]+sumram[44][50]+sumram[44][51]+sumram[44][52]+sumram[44][53]+sumram[44][54]+sumram[44][55]+sumram[44][56]+sumram[44][57]+sumram[44][58]+sumram[44][59]+sumram[44][60]+sumram[44][61]+sumram[44][62]+sumram[44][63]+sumram[44][64]+sumram[44][65]+sumram[44][66]+sumram[44][67]+sumram[44][68]+sumram[44][69]+sumram[44][70]+sumram[44][71]+sumram[44][72]+sumram[44][73]+sumram[44][74]+sumram[44][75]+sumram[44][76]+sumram[44][77]+sumram[44][78]+sumram[44][79]+sumram[44][80]+sumram[44][81]+sumram[44][82]+sumram[44][83]+sumram[44][84]+sumram[44][85]+sumram[44][86]+sumram[44][87]+sumram[44][88]+sumram[44][89]+sumram[44][90]+sumram[44][91]+sumram[44][92]+sumram[44][93]+sumram[44][94]+sumram[44][95]+sumram[44][96]+sumram[44][97]+sumram[44][98]+sumram[44][99]+sumram[44][100]+sumram[44][101]+sumram[44][102]+sumram[44][103]+sumram[44][104]+sumram[44][105]+sumram[44][106]+sumram[44][107]+sumram[44][108]+sumram[44][109]+sumram[44][110]+sumram[44][111]+sumram[44][112]+sumram[44][113]+sumram[44][114]+sumram[44][115]+sumram[44][116]+sumram[44][117]+sumram[44][118]+sumram[44][119]+sumram[44][120]+sumram[44][121]+sumram[44][122]+sumram[44][123]+sumram[44][124]+sumram[44][125]+sumram[44][126]+sumram[44][127]+sumram[44][128]+sumram[44][129]+sumram[44][130]+sumram[44][131]+sumram[44][132]+sumram[44][133]+sumram[44][134]+sumram[44][135]+sumram[44][136];
    assign sumcache[45]=sumram[45][0]+sumram[45][1]+sumram[45][2]+sumram[45][3]+sumram[45][4]+sumram[45][5]+sumram[45][6]+sumram[45][7]+sumram[45][8]+sumram[45][9]+sumram[45][10]+sumram[45][11]+sumram[45][12]+sumram[45][13]+sumram[45][14]+sumram[45][15]+sumram[45][16]+sumram[45][17]+sumram[45][18]+sumram[45][19]+sumram[45][20]+sumram[45][21]+sumram[45][22]+sumram[45][23]+sumram[45][24]+sumram[45][25]+sumram[45][26]+sumram[45][27]+sumram[45][28]+sumram[45][29]+sumram[45][30]+sumram[45][31]+sumram[45][32]+sumram[45][33]+sumram[45][34]+sumram[45][35]+sumram[45][36]+sumram[45][37]+sumram[45][38]+sumram[45][39]+sumram[45][40]+sumram[45][41]+sumram[45][42]+sumram[45][43]+sumram[45][44]+sumram[45][45]+sumram[45][46]+sumram[45][47]+sumram[45][48]+sumram[45][49]+sumram[45][50]+sumram[45][51]+sumram[45][52]+sumram[45][53]+sumram[45][54]+sumram[45][55]+sumram[45][56]+sumram[45][57]+sumram[45][58]+sumram[45][59]+sumram[45][60]+sumram[45][61]+sumram[45][62]+sumram[45][63]+sumram[45][64]+sumram[45][65]+sumram[45][66]+sumram[45][67]+sumram[45][68]+sumram[45][69]+sumram[45][70]+sumram[45][71]+sumram[45][72]+sumram[45][73]+sumram[45][74]+sumram[45][75]+sumram[45][76]+sumram[45][77]+sumram[45][78]+sumram[45][79]+sumram[45][80]+sumram[45][81]+sumram[45][82]+sumram[45][83]+sumram[45][84]+sumram[45][85]+sumram[45][86]+sumram[45][87]+sumram[45][88]+sumram[45][89]+sumram[45][90]+sumram[45][91]+sumram[45][92]+sumram[45][93]+sumram[45][94]+sumram[45][95]+sumram[45][96]+sumram[45][97]+sumram[45][98]+sumram[45][99]+sumram[45][100]+sumram[45][101]+sumram[45][102]+sumram[45][103]+sumram[45][104]+sumram[45][105]+sumram[45][106]+sumram[45][107]+sumram[45][108]+sumram[45][109]+sumram[45][110]+sumram[45][111]+sumram[45][112]+sumram[45][113]+sumram[45][114]+sumram[45][115]+sumram[45][116]+sumram[45][117]+sumram[45][118]+sumram[45][119]+sumram[45][120]+sumram[45][121]+sumram[45][122]+sumram[45][123]+sumram[45][124]+sumram[45][125]+sumram[45][126]+sumram[45][127]+sumram[45][128]+sumram[45][129]+sumram[45][130]+sumram[45][131]+sumram[45][132]+sumram[45][133]+sumram[45][134]+sumram[45][135]+sumram[45][136];
    assign sumcache[46]=sumram[46][0]+sumram[46][1]+sumram[46][2]+sumram[46][3]+sumram[46][4]+sumram[46][5]+sumram[46][6]+sumram[46][7]+sumram[46][8]+sumram[46][9]+sumram[46][10]+sumram[46][11]+sumram[46][12]+sumram[46][13]+sumram[46][14]+sumram[46][15]+sumram[46][16]+sumram[46][17]+sumram[46][18]+sumram[46][19]+sumram[46][20]+sumram[46][21]+sumram[46][22]+sumram[46][23]+sumram[46][24]+sumram[46][25]+sumram[46][26]+sumram[46][27]+sumram[46][28]+sumram[46][29]+sumram[46][30]+sumram[46][31]+sumram[46][32]+sumram[46][33]+sumram[46][34]+sumram[46][35]+sumram[46][36]+sumram[46][37]+sumram[46][38]+sumram[46][39]+sumram[46][40]+sumram[46][41]+sumram[46][42]+sumram[46][43]+sumram[46][44]+sumram[46][45]+sumram[46][46]+sumram[46][47]+sumram[46][48]+sumram[46][49]+sumram[46][50]+sumram[46][51]+sumram[46][52]+sumram[46][53]+sumram[46][54]+sumram[46][55]+sumram[46][56]+sumram[46][57]+sumram[46][58]+sumram[46][59]+sumram[46][60]+sumram[46][61]+sumram[46][62]+sumram[46][63]+sumram[46][64]+sumram[46][65]+sumram[46][66]+sumram[46][67]+sumram[46][68]+sumram[46][69]+sumram[46][70]+sumram[46][71]+sumram[46][72]+sumram[46][73]+sumram[46][74]+sumram[46][75]+sumram[46][76]+sumram[46][77]+sumram[46][78]+sumram[46][79]+sumram[46][80]+sumram[46][81]+sumram[46][82]+sumram[46][83]+sumram[46][84]+sumram[46][85]+sumram[46][86]+sumram[46][87]+sumram[46][88]+sumram[46][89]+sumram[46][90]+sumram[46][91]+sumram[46][92]+sumram[46][93]+sumram[46][94]+sumram[46][95]+sumram[46][96]+sumram[46][97]+sumram[46][98]+sumram[46][99]+sumram[46][100]+sumram[46][101]+sumram[46][102]+sumram[46][103]+sumram[46][104]+sumram[46][105]+sumram[46][106]+sumram[46][107]+sumram[46][108]+sumram[46][109]+sumram[46][110]+sumram[46][111]+sumram[46][112]+sumram[46][113]+sumram[46][114]+sumram[46][115]+sumram[46][116]+sumram[46][117]+sumram[46][118]+sumram[46][119]+sumram[46][120]+sumram[46][121]+sumram[46][122]+sumram[46][123]+sumram[46][124]+sumram[46][125]+sumram[46][126]+sumram[46][127]+sumram[46][128]+sumram[46][129]+sumram[46][130]+sumram[46][131]+sumram[46][132]+sumram[46][133]+sumram[46][134]+sumram[46][135]+sumram[46][136];
    assign sumcache[47]=sumram[47][0]+sumram[47][1]+sumram[47][2]+sumram[47][3]+sumram[47][4]+sumram[47][5]+sumram[47][6]+sumram[47][7]+sumram[47][8]+sumram[47][9]+sumram[47][10]+sumram[47][11]+sumram[47][12]+sumram[47][13]+sumram[47][14]+sumram[47][15]+sumram[47][16]+sumram[47][17]+sumram[47][18]+sumram[47][19]+sumram[47][20]+sumram[47][21]+sumram[47][22]+sumram[47][23]+sumram[47][24]+sumram[47][25]+sumram[47][26]+sumram[47][27]+sumram[47][28]+sumram[47][29]+sumram[47][30]+sumram[47][31]+sumram[47][32]+sumram[47][33]+sumram[47][34]+sumram[47][35]+sumram[47][36]+sumram[47][37]+sumram[47][38]+sumram[47][39]+sumram[47][40]+sumram[47][41]+sumram[47][42]+sumram[47][43]+sumram[47][44]+sumram[47][45]+sumram[47][46]+sumram[47][47]+sumram[47][48]+sumram[47][49]+sumram[47][50]+sumram[47][51]+sumram[47][52]+sumram[47][53]+sumram[47][54]+sumram[47][55]+sumram[47][56]+sumram[47][57]+sumram[47][58]+sumram[47][59]+sumram[47][60]+sumram[47][61]+sumram[47][62]+sumram[47][63]+sumram[47][64]+sumram[47][65]+sumram[47][66]+sumram[47][67]+sumram[47][68]+sumram[47][69]+sumram[47][70]+sumram[47][71]+sumram[47][72]+sumram[47][73]+sumram[47][74]+sumram[47][75]+sumram[47][76]+sumram[47][77]+sumram[47][78]+sumram[47][79]+sumram[47][80]+sumram[47][81]+sumram[47][82]+sumram[47][83]+sumram[47][84]+sumram[47][85]+sumram[47][86]+sumram[47][87]+sumram[47][88]+sumram[47][89]+sumram[47][90]+sumram[47][91]+sumram[47][92]+sumram[47][93]+sumram[47][94]+sumram[47][95]+sumram[47][96]+sumram[47][97]+sumram[47][98]+sumram[47][99]+sumram[47][100]+sumram[47][101]+sumram[47][102]+sumram[47][103]+sumram[47][104]+sumram[47][105]+sumram[47][106]+sumram[47][107]+sumram[47][108]+sumram[47][109]+sumram[47][110]+sumram[47][111]+sumram[47][112]+sumram[47][113]+sumram[47][114]+sumram[47][115]+sumram[47][116]+sumram[47][117]+sumram[47][118]+sumram[47][119]+sumram[47][120]+sumram[47][121]+sumram[47][122]+sumram[47][123]+sumram[47][124]+sumram[47][125]+sumram[47][126]+sumram[47][127]+sumram[47][128]+sumram[47][129]+sumram[47][130]+sumram[47][131]+sumram[47][132]+sumram[47][133]+sumram[47][134]+sumram[47][135]+sumram[47][136];
    assign sumcache[48]=sumram[48][0]+sumram[48][1]+sumram[48][2]+sumram[48][3]+sumram[48][4]+sumram[48][5]+sumram[48][6]+sumram[48][7]+sumram[48][8]+sumram[48][9]+sumram[48][10]+sumram[48][11]+sumram[48][12]+sumram[48][13]+sumram[48][14]+sumram[48][15]+sumram[48][16]+sumram[48][17]+sumram[48][18]+sumram[48][19]+sumram[48][20]+sumram[48][21]+sumram[48][22]+sumram[48][23]+sumram[48][24]+sumram[48][25]+sumram[48][26]+sumram[48][27]+sumram[48][28]+sumram[48][29]+sumram[48][30]+sumram[48][31]+sumram[48][32]+sumram[48][33]+sumram[48][34]+sumram[48][35]+sumram[48][36]+sumram[48][37]+sumram[48][38]+sumram[48][39]+sumram[48][40]+sumram[48][41]+sumram[48][42]+sumram[48][43]+sumram[48][44]+sumram[48][45]+sumram[48][46]+sumram[48][47]+sumram[48][48]+sumram[48][49]+sumram[48][50]+sumram[48][51]+sumram[48][52]+sumram[48][53]+sumram[48][54]+sumram[48][55]+sumram[48][56]+sumram[48][57]+sumram[48][58]+sumram[48][59]+sumram[48][60]+sumram[48][61]+sumram[48][62]+sumram[48][63]+sumram[48][64]+sumram[48][65]+sumram[48][66]+sumram[48][67]+sumram[48][68]+sumram[48][69]+sumram[48][70]+sumram[48][71]+sumram[48][72]+sumram[48][73]+sumram[48][74]+sumram[48][75]+sumram[48][76]+sumram[48][77]+sumram[48][78]+sumram[48][79]+sumram[48][80]+sumram[48][81]+sumram[48][82]+sumram[48][83]+sumram[48][84]+sumram[48][85]+sumram[48][86]+sumram[48][87]+sumram[48][88]+sumram[48][89]+sumram[48][90]+sumram[48][91]+sumram[48][92]+sumram[48][93]+sumram[48][94]+sumram[48][95]+sumram[48][96]+sumram[48][97]+sumram[48][98]+sumram[48][99]+sumram[48][100]+sumram[48][101]+sumram[48][102]+sumram[48][103]+sumram[48][104]+sumram[48][105]+sumram[48][106]+sumram[48][107]+sumram[48][108]+sumram[48][109]+sumram[48][110]+sumram[48][111]+sumram[48][112]+sumram[48][113]+sumram[48][114]+sumram[48][115]+sumram[48][116]+sumram[48][117]+sumram[48][118]+sumram[48][119]+sumram[48][120]+sumram[48][121]+sumram[48][122]+sumram[48][123]+sumram[48][124]+sumram[48][125]+sumram[48][126]+sumram[48][127]+sumram[48][128]+sumram[48][129]+sumram[48][130]+sumram[48][131]+sumram[48][132]+sumram[48][133]+sumram[48][134]+sumram[48][135]+sumram[48][136];
    assign sumcache[49]=sumram[49][0]+sumram[49][1]+sumram[49][2]+sumram[49][3]+sumram[49][4]+sumram[49][5]+sumram[49][6]+sumram[49][7]+sumram[49][8]+sumram[49][9]+sumram[49][10]+sumram[49][11]+sumram[49][12]+sumram[49][13]+sumram[49][14]+sumram[49][15]+sumram[49][16]+sumram[49][17]+sumram[49][18]+sumram[49][19]+sumram[49][20]+sumram[49][21]+sumram[49][22]+sumram[49][23]+sumram[49][24]+sumram[49][25]+sumram[49][26]+sumram[49][27]+sumram[49][28]+sumram[49][29]+sumram[49][30]+sumram[49][31]+sumram[49][32]+sumram[49][33]+sumram[49][34]+sumram[49][35]+sumram[49][36]+sumram[49][37]+sumram[49][38]+sumram[49][39]+sumram[49][40]+sumram[49][41]+sumram[49][42]+sumram[49][43]+sumram[49][44]+sumram[49][45]+sumram[49][46]+sumram[49][47]+sumram[49][48]+sumram[49][49]+sumram[49][50]+sumram[49][51]+sumram[49][52]+sumram[49][53]+sumram[49][54]+sumram[49][55]+sumram[49][56]+sumram[49][57]+sumram[49][58]+sumram[49][59]+sumram[49][60]+sumram[49][61]+sumram[49][62]+sumram[49][63]+sumram[49][64]+sumram[49][65]+sumram[49][66]+sumram[49][67]+sumram[49][68]+sumram[49][69]+sumram[49][70]+sumram[49][71]+sumram[49][72]+sumram[49][73]+sumram[49][74]+sumram[49][75]+sumram[49][76]+sumram[49][77]+sumram[49][78]+sumram[49][79]+sumram[49][80]+sumram[49][81]+sumram[49][82]+sumram[49][83]+sumram[49][84]+sumram[49][85]+sumram[49][86]+sumram[49][87]+sumram[49][88]+sumram[49][89]+sumram[49][90]+sumram[49][91]+sumram[49][92]+sumram[49][93]+sumram[49][94]+sumram[49][95]+sumram[49][96]+sumram[49][97]+sumram[49][98]+sumram[49][99]+sumram[49][100]+sumram[49][101]+sumram[49][102]+sumram[49][103]+sumram[49][104]+sumram[49][105]+sumram[49][106]+sumram[49][107]+sumram[49][108]+sumram[49][109]+sumram[49][110]+sumram[49][111]+sumram[49][112]+sumram[49][113]+sumram[49][114]+sumram[49][115]+sumram[49][116]+sumram[49][117]+sumram[49][118]+sumram[49][119]+sumram[49][120]+sumram[49][121]+sumram[49][122]+sumram[49][123]+sumram[49][124]+sumram[49][125]+sumram[49][126]+sumram[49][127]+sumram[49][128]+sumram[49][129]+sumram[49][130]+sumram[49][131]+sumram[49][132]+sumram[49][133]+sumram[49][134]+sumram[49][135]+sumram[49][136];
    assign sumcache[50]=sumram[50][0]+sumram[50][1]+sumram[50][2]+sumram[50][3]+sumram[50][4]+sumram[50][5]+sumram[50][6]+sumram[50][7]+sumram[50][8]+sumram[50][9]+sumram[50][10]+sumram[50][11]+sumram[50][12]+sumram[50][13]+sumram[50][14]+sumram[50][15]+sumram[50][16]+sumram[50][17]+sumram[50][18]+sumram[50][19]+sumram[50][20]+sumram[50][21]+sumram[50][22]+sumram[50][23]+sumram[50][24]+sumram[50][25]+sumram[50][26]+sumram[50][27]+sumram[50][28]+sumram[50][29]+sumram[50][30]+sumram[50][31]+sumram[50][32]+sumram[50][33]+sumram[50][34]+sumram[50][35]+sumram[50][36]+sumram[50][37]+sumram[50][38]+sumram[50][39]+sumram[50][40]+sumram[50][41]+sumram[50][42]+sumram[50][43]+sumram[50][44]+sumram[50][45]+sumram[50][46]+sumram[50][47]+sumram[50][48]+sumram[50][49]+sumram[50][50]+sumram[50][51]+sumram[50][52]+sumram[50][53]+sumram[50][54]+sumram[50][55]+sumram[50][56]+sumram[50][57]+sumram[50][58]+sumram[50][59]+sumram[50][60]+sumram[50][61]+sumram[50][62]+sumram[50][63]+sumram[50][64]+sumram[50][65]+sumram[50][66]+sumram[50][67]+sumram[50][68]+sumram[50][69]+sumram[50][70]+sumram[50][71]+sumram[50][72]+sumram[50][73]+sumram[50][74]+sumram[50][75]+sumram[50][76]+sumram[50][77]+sumram[50][78]+sumram[50][79]+sumram[50][80]+sumram[50][81]+sumram[50][82]+sumram[50][83]+sumram[50][84]+sumram[50][85]+sumram[50][86]+sumram[50][87]+sumram[50][88]+sumram[50][89]+sumram[50][90]+sumram[50][91]+sumram[50][92]+sumram[50][93]+sumram[50][94]+sumram[50][95]+sumram[50][96]+sumram[50][97]+sumram[50][98]+sumram[50][99]+sumram[50][100]+sumram[50][101]+sumram[50][102]+sumram[50][103]+sumram[50][104]+sumram[50][105]+sumram[50][106]+sumram[50][107]+sumram[50][108]+sumram[50][109]+sumram[50][110]+sumram[50][111]+sumram[50][112]+sumram[50][113]+sumram[50][114]+sumram[50][115]+sumram[50][116]+sumram[50][117]+sumram[50][118]+sumram[50][119]+sumram[50][120]+sumram[50][121]+sumram[50][122]+sumram[50][123]+sumram[50][124]+sumram[50][125]+sumram[50][126]+sumram[50][127]+sumram[50][128]+sumram[50][129]+sumram[50][130]+sumram[50][131]+sumram[50][132]+sumram[50][133]+sumram[50][134]+sumram[50][135]+sumram[50][136];
    assign sumcache[51]=sumram[51][0]+sumram[51][1]+sumram[51][2]+sumram[51][3]+sumram[51][4]+sumram[51][5]+sumram[51][6]+sumram[51][7]+sumram[51][8]+sumram[51][9]+sumram[51][10]+sumram[51][11]+sumram[51][12]+sumram[51][13]+sumram[51][14]+sumram[51][15]+sumram[51][16]+sumram[51][17]+sumram[51][18]+sumram[51][19]+sumram[51][20]+sumram[51][21]+sumram[51][22]+sumram[51][23]+sumram[51][24]+sumram[51][25]+sumram[51][26]+sumram[51][27]+sumram[51][28]+sumram[51][29]+sumram[51][30]+sumram[51][31]+sumram[51][32]+sumram[51][33]+sumram[51][34]+sumram[51][35]+sumram[51][36]+sumram[51][37]+sumram[51][38]+sumram[51][39]+sumram[51][40]+sumram[51][41]+sumram[51][42]+sumram[51][43]+sumram[51][44]+sumram[51][45]+sumram[51][46]+sumram[51][47]+sumram[51][48]+sumram[51][49]+sumram[51][50]+sumram[51][51]+sumram[51][52]+sumram[51][53]+sumram[51][54]+sumram[51][55]+sumram[51][56]+sumram[51][57]+sumram[51][58]+sumram[51][59]+sumram[51][60]+sumram[51][61]+sumram[51][62]+sumram[51][63]+sumram[51][64]+sumram[51][65]+sumram[51][66]+sumram[51][67]+sumram[51][68]+sumram[51][69]+sumram[51][70]+sumram[51][71]+sumram[51][72]+sumram[51][73]+sumram[51][74]+sumram[51][75]+sumram[51][76]+sumram[51][77]+sumram[51][78]+sumram[51][79]+sumram[51][80]+sumram[51][81]+sumram[51][82]+sumram[51][83]+sumram[51][84]+sumram[51][85]+sumram[51][86]+sumram[51][87]+sumram[51][88]+sumram[51][89]+sumram[51][90]+sumram[51][91]+sumram[51][92]+sumram[51][93]+sumram[51][94]+sumram[51][95]+sumram[51][96]+sumram[51][97]+sumram[51][98]+sumram[51][99]+sumram[51][100]+sumram[51][101]+sumram[51][102]+sumram[51][103]+sumram[51][104]+sumram[51][105]+sumram[51][106]+sumram[51][107]+sumram[51][108]+sumram[51][109]+sumram[51][110]+sumram[51][111]+sumram[51][112]+sumram[51][113]+sumram[51][114]+sumram[51][115]+sumram[51][116]+sumram[51][117]+sumram[51][118]+sumram[51][119]+sumram[51][120]+sumram[51][121]+sumram[51][122]+sumram[51][123]+sumram[51][124]+sumram[51][125]+sumram[51][126]+sumram[51][127]+sumram[51][128]+sumram[51][129]+sumram[51][130]+sumram[51][131]+sumram[51][132]+sumram[51][133]+sumram[51][134]+sumram[51][135]+sumram[51][136];
    assign sumcache[52]=sumram[52][0]+sumram[52][1]+sumram[52][2]+sumram[52][3]+sumram[52][4]+sumram[52][5]+sumram[52][6]+sumram[52][7]+sumram[52][8]+sumram[52][9]+sumram[52][10]+sumram[52][11]+sumram[52][12]+sumram[52][13]+sumram[52][14]+sumram[52][15]+sumram[52][16]+sumram[52][17]+sumram[52][18]+sumram[52][19]+sumram[52][20]+sumram[52][21]+sumram[52][22]+sumram[52][23]+sumram[52][24]+sumram[52][25]+sumram[52][26]+sumram[52][27]+sumram[52][28]+sumram[52][29]+sumram[52][30]+sumram[52][31]+sumram[52][32]+sumram[52][33]+sumram[52][34]+sumram[52][35]+sumram[52][36]+sumram[52][37]+sumram[52][38]+sumram[52][39]+sumram[52][40]+sumram[52][41]+sumram[52][42]+sumram[52][43]+sumram[52][44]+sumram[52][45]+sumram[52][46]+sumram[52][47]+sumram[52][48]+sumram[52][49]+sumram[52][50]+sumram[52][51]+sumram[52][52]+sumram[52][53]+sumram[52][54]+sumram[52][55]+sumram[52][56]+sumram[52][57]+sumram[52][58]+sumram[52][59]+sumram[52][60]+sumram[52][61]+sumram[52][62]+sumram[52][63]+sumram[52][64]+sumram[52][65]+sumram[52][66]+sumram[52][67]+sumram[52][68]+sumram[52][69]+sumram[52][70]+sumram[52][71]+sumram[52][72]+sumram[52][73]+sumram[52][74]+sumram[52][75]+sumram[52][76]+sumram[52][77]+sumram[52][78]+sumram[52][79]+sumram[52][80]+sumram[52][81]+sumram[52][82]+sumram[52][83]+sumram[52][84]+sumram[52][85]+sumram[52][86]+sumram[52][87]+sumram[52][88]+sumram[52][89]+sumram[52][90]+sumram[52][91]+sumram[52][92]+sumram[52][93]+sumram[52][94]+sumram[52][95]+sumram[52][96]+sumram[52][97]+sumram[52][98]+sumram[52][99]+sumram[52][100]+sumram[52][101]+sumram[52][102]+sumram[52][103]+sumram[52][104]+sumram[52][105]+sumram[52][106]+sumram[52][107]+sumram[52][108]+sumram[52][109]+sumram[52][110]+sumram[52][111]+sumram[52][112]+sumram[52][113]+sumram[52][114]+sumram[52][115]+sumram[52][116]+sumram[52][117]+sumram[52][118]+sumram[52][119]+sumram[52][120]+sumram[52][121]+sumram[52][122]+sumram[52][123]+sumram[52][124]+sumram[52][125]+sumram[52][126]+sumram[52][127]+sumram[52][128]+sumram[52][129]+sumram[52][130]+sumram[52][131]+sumram[52][132]+sumram[52][133]+sumram[52][134]+sumram[52][135]+sumram[52][136];
    assign sumcache[53]=sumram[53][0]+sumram[53][1]+sumram[53][2]+sumram[53][3]+sumram[53][4]+sumram[53][5]+sumram[53][6]+sumram[53][7]+sumram[53][8]+sumram[53][9]+sumram[53][10]+sumram[53][11]+sumram[53][12]+sumram[53][13]+sumram[53][14]+sumram[53][15]+sumram[53][16]+sumram[53][17]+sumram[53][18]+sumram[53][19]+sumram[53][20]+sumram[53][21]+sumram[53][22]+sumram[53][23]+sumram[53][24]+sumram[53][25]+sumram[53][26]+sumram[53][27]+sumram[53][28]+sumram[53][29]+sumram[53][30]+sumram[53][31]+sumram[53][32]+sumram[53][33]+sumram[53][34]+sumram[53][35]+sumram[53][36]+sumram[53][37]+sumram[53][38]+sumram[53][39]+sumram[53][40]+sumram[53][41]+sumram[53][42]+sumram[53][43]+sumram[53][44]+sumram[53][45]+sumram[53][46]+sumram[53][47]+sumram[53][48]+sumram[53][49]+sumram[53][50]+sumram[53][51]+sumram[53][52]+sumram[53][53]+sumram[53][54]+sumram[53][55]+sumram[53][56]+sumram[53][57]+sumram[53][58]+sumram[53][59]+sumram[53][60]+sumram[53][61]+sumram[53][62]+sumram[53][63]+sumram[53][64]+sumram[53][65]+sumram[53][66]+sumram[53][67]+sumram[53][68]+sumram[53][69]+sumram[53][70]+sumram[53][71]+sumram[53][72]+sumram[53][73]+sumram[53][74]+sumram[53][75]+sumram[53][76]+sumram[53][77]+sumram[53][78]+sumram[53][79]+sumram[53][80]+sumram[53][81]+sumram[53][82]+sumram[53][83]+sumram[53][84]+sumram[53][85]+sumram[53][86]+sumram[53][87]+sumram[53][88]+sumram[53][89]+sumram[53][90]+sumram[53][91]+sumram[53][92]+sumram[53][93]+sumram[53][94]+sumram[53][95]+sumram[53][96]+sumram[53][97]+sumram[53][98]+sumram[53][99]+sumram[53][100]+sumram[53][101]+sumram[53][102]+sumram[53][103]+sumram[53][104]+sumram[53][105]+sumram[53][106]+sumram[53][107]+sumram[53][108]+sumram[53][109]+sumram[53][110]+sumram[53][111]+sumram[53][112]+sumram[53][113]+sumram[53][114]+sumram[53][115]+sumram[53][116]+sumram[53][117]+sumram[53][118]+sumram[53][119]+sumram[53][120]+sumram[53][121]+sumram[53][122]+sumram[53][123]+sumram[53][124]+sumram[53][125]+sumram[53][126]+sumram[53][127]+sumram[53][128]+sumram[53][129]+sumram[53][130]+sumram[53][131]+sumram[53][132]+sumram[53][133]+sumram[53][134]+sumram[53][135]+sumram[53][136];
    assign sumcache[54]=sumram[54][0]+sumram[54][1]+sumram[54][2]+sumram[54][3]+sumram[54][4]+sumram[54][5]+sumram[54][6]+sumram[54][7]+sumram[54][8]+sumram[54][9]+sumram[54][10]+sumram[54][11]+sumram[54][12]+sumram[54][13]+sumram[54][14]+sumram[54][15]+sumram[54][16]+sumram[54][17]+sumram[54][18]+sumram[54][19]+sumram[54][20]+sumram[54][21]+sumram[54][22]+sumram[54][23]+sumram[54][24]+sumram[54][25]+sumram[54][26]+sumram[54][27]+sumram[54][28]+sumram[54][29]+sumram[54][30]+sumram[54][31]+sumram[54][32]+sumram[54][33]+sumram[54][34]+sumram[54][35]+sumram[54][36]+sumram[54][37]+sumram[54][38]+sumram[54][39]+sumram[54][40]+sumram[54][41]+sumram[54][42]+sumram[54][43]+sumram[54][44]+sumram[54][45]+sumram[54][46]+sumram[54][47]+sumram[54][48]+sumram[54][49]+sumram[54][50]+sumram[54][51]+sumram[54][52]+sumram[54][53]+sumram[54][54]+sumram[54][55]+sumram[54][56]+sumram[54][57]+sumram[54][58]+sumram[54][59]+sumram[54][60]+sumram[54][61]+sumram[54][62]+sumram[54][63]+sumram[54][64]+sumram[54][65]+sumram[54][66]+sumram[54][67]+sumram[54][68]+sumram[54][69]+sumram[54][70]+sumram[54][71]+sumram[54][72]+sumram[54][73]+sumram[54][74]+sumram[54][75]+sumram[54][76]+sumram[54][77]+sumram[54][78]+sumram[54][79]+sumram[54][80]+sumram[54][81]+sumram[54][82]+sumram[54][83]+sumram[54][84]+sumram[54][85]+sumram[54][86]+sumram[54][87]+sumram[54][88]+sumram[54][89]+sumram[54][90]+sumram[54][91]+sumram[54][92]+sumram[54][93]+sumram[54][94]+sumram[54][95]+sumram[54][96]+sumram[54][97]+sumram[54][98]+sumram[54][99]+sumram[54][100]+sumram[54][101]+sumram[54][102]+sumram[54][103]+sumram[54][104]+sumram[54][105]+sumram[54][106]+sumram[54][107]+sumram[54][108]+sumram[54][109]+sumram[54][110]+sumram[54][111]+sumram[54][112]+sumram[54][113]+sumram[54][114]+sumram[54][115]+sumram[54][116]+sumram[54][117]+sumram[54][118]+sumram[54][119]+sumram[54][120]+sumram[54][121]+sumram[54][122]+sumram[54][123]+sumram[54][124]+sumram[54][125]+sumram[54][126]+sumram[54][127]+sumram[54][128]+sumram[54][129]+sumram[54][130]+sumram[54][131]+sumram[54][132]+sumram[54][133]+sumram[54][134]+sumram[54][135]+sumram[54][136];
    assign sumcache[55]=sumram[55][0]+sumram[55][1]+sumram[55][2]+sumram[55][3]+sumram[55][4]+sumram[55][5]+sumram[55][6]+sumram[55][7]+sumram[55][8]+sumram[55][9]+sumram[55][10]+sumram[55][11]+sumram[55][12]+sumram[55][13]+sumram[55][14]+sumram[55][15]+sumram[55][16]+sumram[55][17]+sumram[55][18]+sumram[55][19]+sumram[55][20]+sumram[55][21]+sumram[55][22]+sumram[55][23]+sumram[55][24]+sumram[55][25]+sumram[55][26]+sumram[55][27]+sumram[55][28]+sumram[55][29]+sumram[55][30]+sumram[55][31]+sumram[55][32]+sumram[55][33]+sumram[55][34]+sumram[55][35]+sumram[55][36]+sumram[55][37]+sumram[55][38]+sumram[55][39]+sumram[55][40]+sumram[55][41]+sumram[55][42]+sumram[55][43]+sumram[55][44]+sumram[55][45]+sumram[55][46]+sumram[55][47]+sumram[55][48]+sumram[55][49]+sumram[55][50]+sumram[55][51]+sumram[55][52]+sumram[55][53]+sumram[55][54]+sumram[55][55]+sumram[55][56]+sumram[55][57]+sumram[55][58]+sumram[55][59]+sumram[55][60]+sumram[55][61]+sumram[55][62]+sumram[55][63]+sumram[55][64]+sumram[55][65]+sumram[55][66]+sumram[55][67]+sumram[55][68]+sumram[55][69]+sumram[55][70]+sumram[55][71]+sumram[55][72]+sumram[55][73]+sumram[55][74]+sumram[55][75]+sumram[55][76]+sumram[55][77]+sumram[55][78]+sumram[55][79]+sumram[55][80]+sumram[55][81]+sumram[55][82]+sumram[55][83]+sumram[55][84]+sumram[55][85]+sumram[55][86]+sumram[55][87]+sumram[55][88]+sumram[55][89]+sumram[55][90]+sumram[55][91]+sumram[55][92]+sumram[55][93]+sumram[55][94]+sumram[55][95]+sumram[55][96]+sumram[55][97]+sumram[55][98]+sumram[55][99]+sumram[55][100]+sumram[55][101]+sumram[55][102]+sumram[55][103]+sumram[55][104]+sumram[55][105]+sumram[55][106]+sumram[55][107]+sumram[55][108]+sumram[55][109]+sumram[55][110]+sumram[55][111]+sumram[55][112]+sumram[55][113]+sumram[55][114]+sumram[55][115]+sumram[55][116]+sumram[55][117]+sumram[55][118]+sumram[55][119]+sumram[55][120]+sumram[55][121]+sumram[55][122]+sumram[55][123]+sumram[55][124]+sumram[55][125]+sumram[55][126]+sumram[55][127]+sumram[55][128]+sumram[55][129]+sumram[55][130]+sumram[55][131]+sumram[55][132]+sumram[55][133]+sumram[55][134]+sumram[55][135]+sumram[55][136];
    assign sumcache[56]=sumram[56][0]+sumram[56][1]+sumram[56][2]+sumram[56][3]+sumram[56][4]+sumram[56][5]+sumram[56][6]+sumram[56][7]+sumram[56][8]+sumram[56][9]+sumram[56][10]+sumram[56][11]+sumram[56][12]+sumram[56][13]+sumram[56][14]+sumram[56][15]+sumram[56][16]+sumram[56][17]+sumram[56][18]+sumram[56][19]+sumram[56][20]+sumram[56][21]+sumram[56][22]+sumram[56][23]+sumram[56][24]+sumram[56][25]+sumram[56][26]+sumram[56][27]+sumram[56][28]+sumram[56][29]+sumram[56][30]+sumram[56][31]+sumram[56][32]+sumram[56][33]+sumram[56][34]+sumram[56][35]+sumram[56][36]+sumram[56][37]+sumram[56][38]+sumram[56][39]+sumram[56][40]+sumram[56][41]+sumram[56][42]+sumram[56][43]+sumram[56][44]+sumram[56][45]+sumram[56][46]+sumram[56][47]+sumram[56][48]+sumram[56][49]+sumram[56][50]+sumram[56][51]+sumram[56][52]+sumram[56][53]+sumram[56][54]+sumram[56][55]+sumram[56][56]+sumram[56][57]+sumram[56][58]+sumram[56][59]+sumram[56][60]+sumram[56][61]+sumram[56][62]+sumram[56][63]+sumram[56][64]+sumram[56][65]+sumram[56][66]+sumram[56][67]+sumram[56][68]+sumram[56][69]+sumram[56][70]+sumram[56][71]+sumram[56][72]+sumram[56][73]+sumram[56][74]+sumram[56][75]+sumram[56][76]+sumram[56][77]+sumram[56][78]+sumram[56][79]+sumram[56][80]+sumram[56][81]+sumram[56][82]+sumram[56][83]+sumram[56][84]+sumram[56][85]+sumram[56][86]+sumram[56][87]+sumram[56][88]+sumram[56][89]+sumram[56][90]+sumram[56][91]+sumram[56][92]+sumram[56][93]+sumram[56][94]+sumram[56][95]+sumram[56][96]+sumram[56][97]+sumram[56][98]+sumram[56][99]+sumram[56][100]+sumram[56][101]+sumram[56][102]+sumram[56][103]+sumram[56][104]+sumram[56][105]+sumram[56][106]+sumram[56][107]+sumram[56][108]+sumram[56][109]+sumram[56][110]+sumram[56][111]+sumram[56][112]+sumram[56][113]+sumram[56][114]+sumram[56][115]+sumram[56][116]+sumram[56][117]+sumram[56][118]+sumram[56][119]+sumram[56][120]+sumram[56][121]+sumram[56][122]+sumram[56][123]+sumram[56][124]+sumram[56][125]+sumram[56][126]+sumram[56][127]+sumram[56][128]+sumram[56][129]+sumram[56][130]+sumram[56][131]+sumram[56][132]+sumram[56][133]+sumram[56][134]+sumram[56][135]+sumram[56][136];
    assign sumcache[57]=sumram[57][0]+sumram[57][1]+sumram[57][2]+sumram[57][3]+sumram[57][4]+sumram[57][5]+sumram[57][6]+sumram[57][7]+sumram[57][8]+sumram[57][9]+sumram[57][10]+sumram[57][11]+sumram[57][12]+sumram[57][13]+sumram[57][14]+sumram[57][15]+sumram[57][16]+sumram[57][17]+sumram[57][18]+sumram[57][19]+sumram[57][20]+sumram[57][21]+sumram[57][22]+sumram[57][23]+sumram[57][24]+sumram[57][25]+sumram[57][26]+sumram[57][27]+sumram[57][28]+sumram[57][29]+sumram[57][30]+sumram[57][31]+sumram[57][32]+sumram[57][33]+sumram[57][34]+sumram[57][35]+sumram[57][36]+sumram[57][37]+sumram[57][38]+sumram[57][39]+sumram[57][40]+sumram[57][41]+sumram[57][42]+sumram[57][43]+sumram[57][44]+sumram[57][45]+sumram[57][46]+sumram[57][47]+sumram[57][48]+sumram[57][49]+sumram[57][50]+sumram[57][51]+sumram[57][52]+sumram[57][53]+sumram[57][54]+sumram[57][55]+sumram[57][56]+sumram[57][57]+sumram[57][58]+sumram[57][59]+sumram[57][60]+sumram[57][61]+sumram[57][62]+sumram[57][63]+sumram[57][64]+sumram[57][65]+sumram[57][66]+sumram[57][67]+sumram[57][68]+sumram[57][69]+sumram[57][70]+sumram[57][71]+sumram[57][72]+sumram[57][73]+sumram[57][74]+sumram[57][75]+sumram[57][76]+sumram[57][77]+sumram[57][78]+sumram[57][79]+sumram[57][80]+sumram[57][81]+sumram[57][82]+sumram[57][83]+sumram[57][84]+sumram[57][85]+sumram[57][86]+sumram[57][87]+sumram[57][88]+sumram[57][89]+sumram[57][90]+sumram[57][91]+sumram[57][92]+sumram[57][93]+sumram[57][94]+sumram[57][95]+sumram[57][96]+sumram[57][97]+sumram[57][98]+sumram[57][99]+sumram[57][100]+sumram[57][101]+sumram[57][102]+sumram[57][103]+sumram[57][104]+sumram[57][105]+sumram[57][106]+sumram[57][107]+sumram[57][108]+sumram[57][109]+sumram[57][110]+sumram[57][111]+sumram[57][112]+sumram[57][113]+sumram[57][114]+sumram[57][115]+sumram[57][116]+sumram[57][117]+sumram[57][118]+sumram[57][119]+sumram[57][120]+sumram[57][121]+sumram[57][122]+sumram[57][123]+sumram[57][124]+sumram[57][125]+sumram[57][126]+sumram[57][127]+sumram[57][128]+sumram[57][129]+sumram[57][130]+sumram[57][131]+sumram[57][132]+sumram[57][133]+sumram[57][134]+sumram[57][135]+sumram[57][136];
    assign sumcache[58]=sumram[58][0]+sumram[58][1]+sumram[58][2]+sumram[58][3]+sumram[58][4]+sumram[58][5]+sumram[58][6]+sumram[58][7]+sumram[58][8]+sumram[58][9]+sumram[58][10]+sumram[58][11]+sumram[58][12]+sumram[58][13]+sumram[58][14]+sumram[58][15]+sumram[58][16]+sumram[58][17]+sumram[58][18]+sumram[58][19]+sumram[58][20]+sumram[58][21]+sumram[58][22]+sumram[58][23]+sumram[58][24]+sumram[58][25]+sumram[58][26]+sumram[58][27]+sumram[58][28]+sumram[58][29]+sumram[58][30]+sumram[58][31]+sumram[58][32]+sumram[58][33]+sumram[58][34]+sumram[58][35]+sumram[58][36]+sumram[58][37]+sumram[58][38]+sumram[58][39]+sumram[58][40]+sumram[58][41]+sumram[58][42]+sumram[58][43]+sumram[58][44]+sumram[58][45]+sumram[58][46]+sumram[58][47]+sumram[58][48]+sumram[58][49]+sumram[58][50]+sumram[58][51]+sumram[58][52]+sumram[58][53]+sumram[58][54]+sumram[58][55]+sumram[58][56]+sumram[58][57]+sumram[58][58]+sumram[58][59]+sumram[58][60]+sumram[58][61]+sumram[58][62]+sumram[58][63]+sumram[58][64]+sumram[58][65]+sumram[58][66]+sumram[58][67]+sumram[58][68]+sumram[58][69]+sumram[58][70]+sumram[58][71]+sumram[58][72]+sumram[58][73]+sumram[58][74]+sumram[58][75]+sumram[58][76]+sumram[58][77]+sumram[58][78]+sumram[58][79]+sumram[58][80]+sumram[58][81]+sumram[58][82]+sumram[58][83]+sumram[58][84]+sumram[58][85]+sumram[58][86]+sumram[58][87]+sumram[58][88]+sumram[58][89]+sumram[58][90]+sumram[58][91]+sumram[58][92]+sumram[58][93]+sumram[58][94]+sumram[58][95]+sumram[58][96]+sumram[58][97]+sumram[58][98]+sumram[58][99]+sumram[58][100]+sumram[58][101]+sumram[58][102]+sumram[58][103]+sumram[58][104]+sumram[58][105]+sumram[58][106]+sumram[58][107]+sumram[58][108]+sumram[58][109]+sumram[58][110]+sumram[58][111]+sumram[58][112]+sumram[58][113]+sumram[58][114]+sumram[58][115]+sumram[58][116]+sumram[58][117]+sumram[58][118]+sumram[58][119]+sumram[58][120]+sumram[58][121]+sumram[58][122]+sumram[58][123]+sumram[58][124]+sumram[58][125]+sumram[58][126]+sumram[58][127]+sumram[58][128]+sumram[58][129]+sumram[58][130]+sumram[58][131]+sumram[58][132]+sumram[58][133]+sumram[58][134]+sumram[58][135]+sumram[58][136];
    assign sumcache[59]=sumram[59][0]+sumram[59][1]+sumram[59][2]+sumram[59][3]+sumram[59][4]+sumram[59][5]+sumram[59][6]+sumram[59][7]+sumram[59][8]+sumram[59][9]+sumram[59][10]+sumram[59][11]+sumram[59][12]+sumram[59][13]+sumram[59][14]+sumram[59][15]+sumram[59][16]+sumram[59][17]+sumram[59][18]+sumram[59][19]+sumram[59][20]+sumram[59][21]+sumram[59][22]+sumram[59][23]+sumram[59][24]+sumram[59][25]+sumram[59][26]+sumram[59][27]+sumram[59][28]+sumram[59][29]+sumram[59][30]+sumram[59][31]+sumram[59][32]+sumram[59][33]+sumram[59][34]+sumram[59][35]+sumram[59][36]+sumram[59][37]+sumram[59][38]+sumram[59][39]+sumram[59][40]+sumram[59][41]+sumram[59][42]+sumram[59][43]+sumram[59][44]+sumram[59][45]+sumram[59][46]+sumram[59][47]+sumram[59][48]+sumram[59][49]+sumram[59][50]+sumram[59][51]+sumram[59][52]+sumram[59][53]+sumram[59][54]+sumram[59][55]+sumram[59][56]+sumram[59][57]+sumram[59][58]+sumram[59][59]+sumram[59][60]+sumram[59][61]+sumram[59][62]+sumram[59][63]+sumram[59][64]+sumram[59][65]+sumram[59][66]+sumram[59][67]+sumram[59][68]+sumram[59][69]+sumram[59][70]+sumram[59][71]+sumram[59][72]+sumram[59][73]+sumram[59][74]+sumram[59][75]+sumram[59][76]+sumram[59][77]+sumram[59][78]+sumram[59][79]+sumram[59][80]+sumram[59][81]+sumram[59][82]+sumram[59][83]+sumram[59][84]+sumram[59][85]+sumram[59][86]+sumram[59][87]+sumram[59][88]+sumram[59][89]+sumram[59][90]+sumram[59][91]+sumram[59][92]+sumram[59][93]+sumram[59][94]+sumram[59][95]+sumram[59][96]+sumram[59][97]+sumram[59][98]+sumram[59][99]+sumram[59][100]+sumram[59][101]+sumram[59][102]+sumram[59][103]+sumram[59][104]+sumram[59][105]+sumram[59][106]+sumram[59][107]+sumram[59][108]+sumram[59][109]+sumram[59][110]+sumram[59][111]+sumram[59][112]+sumram[59][113]+sumram[59][114]+sumram[59][115]+sumram[59][116]+sumram[59][117]+sumram[59][118]+sumram[59][119]+sumram[59][120]+sumram[59][121]+sumram[59][122]+sumram[59][123]+sumram[59][124]+sumram[59][125]+sumram[59][126]+sumram[59][127]+sumram[59][128]+sumram[59][129]+sumram[59][130]+sumram[59][131]+sumram[59][132]+sumram[59][133]+sumram[59][134]+sumram[59][135]+sumram[59][136];
    assign sumcache[60]=sumram[60][0]+sumram[60][1]+sumram[60][2]+sumram[60][3]+sumram[60][4]+sumram[60][5]+sumram[60][6]+sumram[60][7]+sumram[60][8]+sumram[60][9]+sumram[60][10]+sumram[60][11]+sumram[60][12]+sumram[60][13]+sumram[60][14]+sumram[60][15]+sumram[60][16]+sumram[60][17]+sumram[60][18]+sumram[60][19]+sumram[60][20]+sumram[60][21]+sumram[60][22]+sumram[60][23]+sumram[60][24]+sumram[60][25]+sumram[60][26]+sumram[60][27]+sumram[60][28]+sumram[60][29]+sumram[60][30]+sumram[60][31]+sumram[60][32]+sumram[60][33]+sumram[60][34]+sumram[60][35]+sumram[60][36]+sumram[60][37]+sumram[60][38]+sumram[60][39]+sumram[60][40]+sumram[60][41]+sumram[60][42]+sumram[60][43]+sumram[60][44]+sumram[60][45]+sumram[60][46]+sumram[60][47]+sumram[60][48]+sumram[60][49]+sumram[60][50]+sumram[60][51]+sumram[60][52]+sumram[60][53]+sumram[60][54]+sumram[60][55]+sumram[60][56]+sumram[60][57]+sumram[60][58]+sumram[60][59]+sumram[60][60]+sumram[60][61]+sumram[60][62]+sumram[60][63]+sumram[60][64]+sumram[60][65]+sumram[60][66]+sumram[60][67]+sumram[60][68]+sumram[60][69]+sumram[60][70]+sumram[60][71]+sumram[60][72]+sumram[60][73]+sumram[60][74]+sumram[60][75]+sumram[60][76]+sumram[60][77]+sumram[60][78]+sumram[60][79]+sumram[60][80]+sumram[60][81]+sumram[60][82]+sumram[60][83]+sumram[60][84]+sumram[60][85]+sumram[60][86]+sumram[60][87]+sumram[60][88]+sumram[60][89]+sumram[60][90]+sumram[60][91]+sumram[60][92]+sumram[60][93]+sumram[60][94]+sumram[60][95]+sumram[60][96]+sumram[60][97]+sumram[60][98]+sumram[60][99]+sumram[60][100]+sumram[60][101]+sumram[60][102]+sumram[60][103]+sumram[60][104]+sumram[60][105]+sumram[60][106]+sumram[60][107]+sumram[60][108]+sumram[60][109]+sumram[60][110]+sumram[60][111]+sumram[60][112]+sumram[60][113]+sumram[60][114]+sumram[60][115]+sumram[60][116]+sumram[60][117]+sumram[60][118]+sumram[60][119]+sumram[60][120]+sumram[60][121]+sumram[60][122]+sumram[60][123]+sumram[60][124]+sumram[60][125]+sumram[60][126]+sumram[60][127]+sumram[60][128]+sumram[60][129]+sumram[60][130]+sumram[60][131]+sumram[60][132]+sumram[60][133]+sumram[60][134]+sumram[60][135]+sumram[60][136];
    assign sumcache[61]=sumram[61][0]+sumram[61][1]+sumram[61][2]+sumram[61][3]+sumram[61][4]+sumram[61][5]+sumram[61][6]+sumram[61][7]+sumram[61][8]+sumram[61][9]+sumram[61][10]+sumram[61][11]+sumram[61][12]+sumram[61][13]+sumram[61][14]+sumram[61][15]+sumram[61][16]+sumram[61][17]+sumram[61][18]+sumram[61][19]+sumram[61][20]+sumram[61][21]+sumram[61][22]+sumram[61][23]+sumram[61][24]+sumram[61][25]+sumram[61][26]+sumram[61][27]+sumram[61][28]+sumram[61][29]+sumram[61][30]+sumram[61][31]+sumram[61][32]+sumram[61][33]+sumram[61][34]+sumram[61][35]+sumram[61][36]+sumram[61][37]+sumram[61][38]+sumram[61][39]+sumram[61][40]+sumram[61][41]+sumram[61][42]+sumram[61][43]+sumram[61][44]+sumram[61][45]+sumram[61][46]+sumram[61][47]+sumram[61][48]+sumram[61][49]+sumram[61][50]+sumram[61][51]+sumram[61][52]+sumram[61][53]+sumram[61][54]+sumram[61][55]+sumram[61][56]+sumram[61][57]+sumram[61][58]+sumram[61][59]+sumram[61][60]+sumram[61][61]+sumram[61][62]+sumram[61][63]+sumram[61][64]+sumram[61][65]+sumram[61][66]+sumram[61][67]+sumram[61][68]+sumram[61][69]+sumram[61][70]+sumram[61][71]+sumram[61][72]+sumram[61][73]+sumram[61][74]+sumram[61][75]+sumram[61][76]+sumram[61][77]+sumram[61][78]+sumram[61][79]+sumram[61][80]+sumram[61][81]+sumram[61][82]+sumram[61][83]+sumram[61][84]+sumram[61][85]+sumram[61][86]+sumram[61][87]+sumram[61][88]+sumram[61][89]+sumram[61][90]+sumram[61][91]+sumram[61][92]+sumram[61][93]+sumram[61][94]+sumram[61][95]+sumram[61][96]+sumram[61][97]+sumram[61][98]+sumram[61][99]+sumram[61][100]+sumram[61][101]+sumram[61][102]+sumram[61][103]+sumram[61][104]+sumram[61][105]+sumram[61][106]+sumram[61][107]+sumram[61][108]+sumram[61][109]+sumram[61][110]+sumram[61][111]+sumram[61][112]+sumram[61][113]+sumram[61][114]+sumram[61][115]+sumram[61][116]+sumram[61][117]+sumram[61][118]+sumram[61][119]+sumram[61][120]+sumram[61][121]+sumram[61][122]+sumram[61][123]+sumram[61][124]+sumram[61][125]+sumram[61][126]+sumram[61][127]+sumram[61][128]+sumram[61][129]+sumram[61][130]+sumram[61][131]+sumram[61][132]+sumram[61][133]+sumram[61][134]+sumram[61][135]+sumram[61][136];
    assign sumcache[62]=sumram[62][0]+sumram[62][1]+sumram[62][2]+sumram[62][3]+sumram[62][4]+sumram[62][5]+sumram[62][6]+sumram[62][7]+sumram[62][8]+sumram[62][9]+sumram[62][10]+sumram[62][11]+sumram[62][12]+sumram[62][13]+sumram[62][14]+sumram[62][15]+sumram[62][16]+sumram[62][17]+sumram[62][18]+sumram[62][19]+sumram[62][20]+sumram[62][21]+sumram[62][22]+sumram[62][23]+sumram[62][24]+sumram[62][25]+sumram[62][26]+sumram[62][27]+sumram[62][28]+sumram[62][29]+sumram[62][30]+sumram[62][31]+sumram[62][32]+sumram[62][33]+sumram[62][34]+sumram[62][35]+sumram[62][36]+sumram[62][37]+sumram[62][38]+sumram[62][39]+sumram[62][40]+sumram[62][41]+sumram[62][42]+sumram[62][43]+sumram[62][44]+sumram[62][45]+sumram[62][46]+sumram[62][47]+sumram[62][48]+sumram[62][49]+sumram[62][50]+sumram[62][51]+sumram[62][52]+sumram[62][53]+sumram[62][54]+sumram[62][55]+sumram[62][56]+sumram[62][57]+sumram[62][58]+sumram[62][59]+sumram[62][60]+sumram[62][61]+sumram[62][62]+sumram[62][63]+sumram[62][64]+sumram[62][65]+sumram[62][66]+sumram[62][67]+sumram[62][68]+sumram[62][69]+sumram[62][70]+sumram[62][71]+sumram[62][72]+sumram[62][73]+sumram[62][74]+sumram[62][75]+sumram[62][76]+sumram[62][77]+sumram[62][78]+sumram[62][79]+sumram[62][80]+sumram[62][81]+sumram[62][82]+sumram[62][83]+sumram[62][84]+sumram[62][85]+sumram[62][86]+sumram[62][87]+sumram[62][88]+sumram[62][89]+sumram[62][90]+sumram[62][91]+sumram[62][92]+sumram[62][93]+sumram[62][94]+sumram[62][95]+sumram[62][96]+sumram[62][97]+sumram[62][98]+sumram[62][99]+sumram[62][100]+sumram[62][101]+sumram[62][102]+sumram[62][103]+sumram[62][104]+sumram[62][105]+sumram[62][106]+sumram[62][107]+sumram[62][108]+sumram[62][109]+sumram[62][110]+sumram[62][111]+sumram[62][112]+sumram[62][113]+sumram[62][114]+sumram[62][115]+sumram[62][116]+sumram[62][117]+sumram[62][118]+sumram[62][119]+sumram[62][120]+sumram[62][121]+sumram[62][122]+sumram[62][123]+sumram[62][124]+sumram[62][125]+sumram[62][126]+sumram[62][127]+sumram[62][128]+sumram[62][129]+sumram[62][130]+sumram[62][131]+sumram[62][132]+sumram[62][133]+sumram[62][134]+sumram[62][135]+sumram[62][136];
    assign sumcache[63]=sumram[63][0]+sumram[63][1]+sumram[63][2]+sumram[63][3]+sumram[63][4]+sumram[63][5]+sumram[63][6]+sumram[63][7]+sumram[63][8]+sumram[63][9]+sumram[63][10]+sumram[63][11]+sumram[63][12]+sumram[63][13]+sumram[63][14]+sumram[63][15]+sumram[63][16]+sumram[63][17]+sumram[63][18]+sumram[63][19]+sumram[63][20]+sumram[63][21]+sumram[63][22]+sumram[63][23]+sumram[63][24]+sumram[63][25]+sumram[63][26]+sumram[63][27]+sumram[63][28]+sumram[63][29]+sumram[63][30]+sumram[63][31]+sumram[63][32]+sumram[63][33]+sumram[63][34]+sumram[63][35]+sumram[63][36]+sumram[63][37]+sumram[63][38]+sumram[63][39]+sumram[63][40]+sumram[63][41]+sumram[63][42]+sumram[63][43]+sumram[63][44]+sumram[63][45]+sumram[63][46]+sumram[63][47]+sumram[63][48]+sumram[63][49]+sumram[63][50]+sumram[63][51]+sumram[63][52]+sumram[63][53]+sumram[63][54]+sumram[63][55]+sumram[63][56]+sumram[63][57]+sumram[63][58]+sumram[63][59]+sumram[63][60]+sumram[63][61]+sumram[63][62]+sumram[63][63]+sumram[63][64]+sumram[63][65]+sumram[63][66]+sumram[63][67]+sumram[63][68]+sumram[63][69]+sumram[63][70]+sumram[63][71]+sumram[63][72]+sumram[63][73]+sumram[63][74]+sumram[63][75]+sumram[63][76]+sumram[63][77]+sumram[63][78]+sumram[63][79]+sumram[63][80]+sumram[63][81]+sumram[63][82]+sumram[63][83]+sumram[63][84]+sumram[63][85]+sumram[63][86]+sumram[63][87]+sumram[63][88]+sumram[63][89]+sumram[63][90]+sumram[63][91]+sumram[63][92]+sumram[63][93]+sumram[63][94]+sumram[63][95]+sumram[63][96]+sumram[63][97]+sumram[63][98]+sumram[63][99]+sumram[63][100]+sumram[63][101]+sumram[63][102]+sumram[63][103]+sumram[63][104]+sumram[63][105]+sumram[63][106]+sumram[63][107]+sumram[63][108]+sumram[63][109]+sumram[63][110]+sumram[63][111]+sumram[63][112]+sumram[63][113]+sumram[63][114]+sumram[63][115]+sumram[63][116]+sumram[63][117]+sumram[63][118]+sumram[63][119]+sumram[63][120]+sumram[63][121]+sumram[63][122]+sumram[63][123]+sumram[63][124]+sumram[63][125]+sumram[63][126]+sumram[63][127]+sumram[63][128]+sumram[63][129]+sumram[63][130]+sumram[63][131]+sumram[63][132]+sumram[63][133]+sumram[63][134]+sumram[63][135]+sumram[63][136];
    assign sumcache[64]=sumram[64][0]+sumram[64][1]+sumram[64][2]+sumram[64][3]+sumram[64][4]+sumram[64][5]+sumram[64][6]+sumram[64][7]+sumram[64][8]+sumram[64][9]+sumram[64][10]+sumram[64][11]+sumram[64][12]+sumram[64][13]+sumram[64][14]+sumram[64][15]+sumram[64][16]+sumram[64][17]+sumram[64][18]+sumram[64][19]+sumram[64][20]+sumram[64][21]+sumram[64][22]+sumram[64][23]+sumram[64][24]+sumram[64][25]+sumram[64][26]+sumram[64][27]+sumram[64][28]+sumram[64][29]+sumram[64][30]+sumram[64][31]+sumram[64][32]+sumram[64][33]+sumram[64][34]+sumram[64][35]+sumram[64][36]+sumram[64][37]+sumram[64][38]+sumram[64][39]+sumram[64][40]+sumram[64][41]+sumram[64][42]+sumram[64][43]+sumram[64][44]+sumram[64][45]+sumram[64][46]+sumram[64][47]+sumram[64][48]+sumram[64][49]+sumram[64][50]+sumram[64][51]+sumram[64][52]+sumram[64][53]+sumram[64][54]+sumram[64][55]+sumram[64][56]+sumram[64][57]+sumram[64][58]+sumram[64][59]+sumram[64][60]+sumram[64][61]+sumram[64][62]+sumram[64][63]+sumram[64][64]+sumram[64][65]+sumram[64][66]+sumram[64][67]+sumram[64][68]+sumram[64][69]+sumram[64][70]+sumram[64][71]+sumram[64][72]+sumram[64][73]+sumram[64][74]+sumram[64][75]+sumram[64][76]+sumram[64][77]+sumram[64][78]+sumram[64][79]+sumram[64][80]+sumram[64][81]+sumram[64][82]+sumram[64][83]+sumram[64][84]+sumram[64][85]+sumram[64][86]+sumram[64][87]+sumram[64][88]+sumram[64][89]+sumram[64][90]+sumram[64][91]+sumram[64][92]+sumram[64][93]+sumram[64][94]+sumram[64][95]+sumram[64][96]+sumram[64][97]+sumram[64][98]+sumram[64][99]+sumram[64][100]+sumram[64][101]+sumram[64][102]+sumram[64][103]+sumram[64][104]+sumram[64][105]+sumram[64][106]+sumram[64][107]+sumram[64][108]+sumram[64][109]+sumram[64][110]+sumram[64][111]+sumram[64][112]+sumram[64][113]+sumram[64][114]+sumram[64][115]+sumram[64][116]+sumram[64][117]+sumram[64][118]+sumram[64][119]+sumram[64][120]+sumram[64][121]+sumram[64][122]+sumram[64][123]+sumram[64][124]+sumram[64][125]+sumram[64][126]+sumram[64][127]+sumram[64][128]+sumram[64][129]+sumram[64][130]+sumram[64][131]+sumram[64][132]+sumram[64][133]+sumram[64][134]+sumram[64][135]+sumram[64][136];
    assign sumcache[65]=sumram[65][0]+sumram[65][1]+sumram[65][2]+sumram[65][3]+sumram[65][4]+sumram[65][5]+sumram[65][6]+sumram[65][7]+sumram[65][8]+sumram[65][9]+sumram[65][10]+sumram[65][11]+sumram[65][12]+sumram[65][13]+sumram[65][14]+sumram[65][15]+sumram[65][16]+sumram[65][17]+sumram[65][18]+sumram[65][19]+sumram[65][20]+sumram[65][21]+sumram[65][22]+sumram[65][23]+sumram[65][24]+sumram[65][25]+sumram[65][26]+sumram[65][27]+sumram[65][28]+sumram[65][29]+sumram[65][30]+sumram[65][31]+sumram[65][32]+sumram[65][33]+sumram[65][34]+sumram[65][35]+sumram[65][36]+sumram[65][37]+sumram[65][38]+sumram[65][39]+sumram[65][40]+sumram[65][41]+sumram[65][42]+sumram[65][43]+sumram[65][44]+sumram[65][45]+sumram[65][46]+sumram[65][47]+sumram[65][48]+sumram[65][49]+sumram[65][50]+sumram[65][51]+sumram[65][52]+sumram[65][53]+sumram[65][54]+sumram[65][55]+sumram[65][56]+sumram[65][57]+sumram[65][58]+sumram[65][59]+sumram[65][60]+sumram[65][61]+sumram[65][62]+sumram[65][63]+sumram[65][64]+sumram[65][65]+sumram[65][66]+sumram[65][67]+sumram[65][68]+sumram[65][69]+sumram[65][70]+sumram[65][71]+sumram[65][72]+sumram[65][73]+sumram[65][74]+sumram[65][75]+sumram[65][76]+sumram[65][77]+sumram[65][78]+sumram[65][79]+sumram[65][80]+sumram[65][81]+sumram[65][82]+sumram[65][83]+sumram[65][84]+sumram[65][85]+sumram[65][86]+sumram[65][87]+sumram[65][88]+sumram[65][89]+sumram[65][90]+sumram[65][91]+sumram[65][92]+sumram[65][93]+sumram[65][94]+sumram[65][95]+sumram[65][96]+sumram[65][97]+sumram[65][98]+sumram[65][99]+sumram[65][100]+sumram[65][101]+sumram[65][102]+sumram[65][103]+sumram[65][104]+sumram[65][105]+sumram[65][106]+sumram[65][107]+sumram[65][108]+sumram[65][109]+sumram[65][110]+sumram[65][111]+sumram[65][112]+sumram[65][113]+sumram[65][114]+sumram[65][115]+sumram[65][116]+sumram[65][117]+sumram[65][118]+sumram[65][119]+sumram[65][120]+sumram[65][121]+sumram[65][122]+sumram[65][123]+sumram[65][124]+sumram[65][125]+sumram[65][126]+sumram[65][127]+sumram[65][128]+sumram[65][129]+sumram[65][130]+sumram[65][131]+sumram[65][132]+sumram[65][133]+sumram[65][134]+sumram[65][135]+sumram[65][136];
    assign sumcache[66]=sumram[66][0]+sumram[66][1]+sumram[66][2]+sumram[66][3]+sumram[66][4]+sumram[66][5]+sumram[66][6]+sumram[66][7]+sumram[66][8]+sumram[66][9]+sumram[66][10]+sumram[66][11]+sumram[66][12]+sumram[66][13]+sumram[66][14]+sumram[66][15]+sumram[66][16]+sumram[66][17]+sumram[66][18]+sumram[66][19]+sumram[66][20]+sumram[66][21]+sumram[66][22]+sumram[66][23]+sumram[66][24]+sumram[66][25]+sumram[66][26]+sumram[66][27]+sumram[66][28]+sumram[66][29]+sumram[66][30]+sumram[66][31]+sumram[66][32]+sumram[66][33]+sumram[66][34]+sumram[66][35]+sumram[66][36]+sumram[66][37]+sumram[66][38]+sumram[66][39]+sumram[66][40]+sumram[66][41]+sumram[66][42]+sumram[66][43]+sumram[66][44]+sumram[66][45]+sumram[66][46]+sumram[66][47]+sumram[66][48]+sumram[66][49]+sumram[66][50]+sumram[66][51]+sumram[66][52]+sumram[66][53]+sumram[66][54]+sumram[66][55]+sumram[66][56]+sumram[66][57]+sumram[66][58]+sumram[66][59]+sumram[66][60]+sumram[66][61]+sumram[66][62]+sumram[66][63]+sumram[66][64]+sumram[66][65]+sumram[66][66]+sumram[66][67]+sumram[66][68]+sumram[66][69]+sumram[66][70]+sumram[66][71]+sumram[66][72]+sumram[66][73]+sumram[66][74]+sumram[66][75]+sumram[66][76]+sumram[66][77]+sumram[66][78]+sumram[66][79]+sumram[66][80]+sumram[66][81]+sumram[66][82]+sumram[66][83]+sumram[66][84]+sumram[66][85]+sumram[66][86]+sumram[66][87]+sumram[66][88]+sumram[66][89]+sumram[66][90]+sumram[66][91]+sumram[66][92]+sumram[66][93]+sumram[66][94]+sumram[66][95]+sumram[66][96]+sumram[66][97]+sumram[66][98]+sumram[66][99]+sumram[66][100]+sumram[66][101]+sumram[66][102]+sumram[66][103]+sumram[66][104]+sumram[66][105]+sumram[66][106]+sumram[66][107]+sumram[66][108]+sumram[66][109]+sumram[66][110]+sumram[66][111]+sumram[66][112]+sumram[66][113]+sumram[66][114]+sumram[66][115]+sumram[66][116]+sumram[66][117]+sumram[66][118]+sumram[66][119]+sumram[66][120]+sumram[66][121]+sumram[66][122]+sumram[66][123]+sumram[66][124]+sumram[66][125]+sumram[66][126]+sumram[66][127]+sumram[66][128]+sumram[66][129]+sumram[66][130]+sumram[66][131]+sumram[66][132]+sumram[66][133]+sumram[66][134]+sumram[66][135]+sumram[66][136];
    assign sumcache[67]=sumram[67][0]+sumram[67][1]+sumram[67][2]+sumram[67][3]+sumram[67][4]+sumram[67][5]+sumram[67][6]+sumram[67][7]+sumram[67][8]+sumram[67][9]+sumram[67][10]+sumram[67][11]+sumram[67][12]+sumram[67][13]+sumram[67][14]+sumram[67][15]+sumram[67][16]+sumram[67][17]+sumram[67][18]+sumram[67][19]+sumram[67][20]+sumram[67][21]+sumram[67][22]+sumram[67][23]+sumram[67][24]+sumram[67][25]+sumram[67][26]+sumram[67][27]+sumram[67][28]+sumram[67][29]+sumram[67][30]+sumram[67][31]+sumram[67][32]+sumram[67][33]+sumram[67][34]+sumram[67][35]+sumram[67][36]+sumram[67][37]+sumram[67][38]+sumram[67][39]+sumram[67][40]+sumram[67][41]+sumram[67][42]+sumram[67][43]+sumram[67][44]+sumram[67][45]+sumram[67][46]+sumram[67][47]+sumram[67][48]+sumram[67][49]+sumram[67][50]+sumram[67][51]+sumram[67][52]+sumram[67][53]+sumram[67][54]+sumram[67][55]+sumram[67][56]+sumram[67][57]+sumram[67][58]+sumram[67][59]+sumram[67][60]+sumram[67][61]+sumram[67][62]+sumram[67][63]+sumram[67][64]+sumram[67][65]+sumram[67][66]+sumram[67][67]+sumram[67][68]+sumram[67][69]+sumram[67][70]+sumram[67][71]+sumram[67][72]+sumram[67][73]+sumram[67][74]+sumram[67][75]+sumram[67][76]+sumram[67][77]+sumram[67][78]+sumram[67][79]+sumram[67][80]+sumram[67][81]+sumram[67][82]+sumram[67][83]+sumram[67][84]+sumram[67][85]+sumram[67][86]+sumram[67][87]+sumram[67][88]+sumram[67][89]+sumram[67][90]+sumram[67][91]+sumram[67][92]+sumram[67][93]+sumram[67][94]+sumram[67][95]+sumram[67][96]+sumram[67][97]+sumram[67][98]+sumram[67][99]+sumram[67][100]+sumram[67][101]+sumram[67][102]+sumram[67][103]+sumram[67][104]+sumram[67][105]+sumram[67][106]+sumram[67][107]+sumram[67][108]+sumram[67][109]+sumram[67][110]+sumram[67][111]+sumram[67][112]+sumram[67][113]+sumram[67][114]+sumram[67][115]+sumram[67][116]+sumram[67][117]+sumram[67][118]+sumram[67][119]+sumram[67][120]+sumram[67][121]+sumram[67][122]+sumram[67][123]+sumram[67][124]+sumram[67][125]+sumram[67][126]+sumram[67][127]+sumram[67][128]+sumram[67][129]+sumram[67][130]+sumram[67][131]+sumram[67][132]+sumram[67][133]+sumram[67][134]+sumram[67][135]+sumram[67][136];
    assign sumcache[68]=sumram[68][0]+sumram[68][1]+sumram[68][2]+sumram[68][3]+sumram[68][4]+sumram[68][5]+sumram[68][6]+sumram[68][7]+sumram[68][8]+sumram[68][9]+sumram[68][10]+sumram[68][11]+sumram[68][12]+sumram[68][13]+sumram[68][14]+sumram[68][15]+sumram[68][16]+sumram[68][17]+sumram[68][18]+sumram[68][19]+sumram[68][20]+sumram[68][21]+sumram[68][22]+sumram[68][23]+sumram[68][24]+sumram[68][25]+sumram[68][26]+sumram[68][27]+sumram[68][28]+sumram[68][29]+sumram[68][30]+sumram[68][31]+sumram[68][32]+sumram[68][33]+sumram[68][34]+sumram[68][35]+sumram[68][36]+sumram[68][37]+sumram[68][38]+sumram[68][39]+sumram[68][40]+sumram[68][41]+sumram[68][42]+sumram[68][43]+sumram[68][44]+sumram[68][45]+sumram[68][46]+sumram[68][47]+sumram[68][48]+sumram[68][49]+sumram[68][50]+sumram[68][51]+sumram[68][52]+sumram[68][53]+sumram[68][54]+sumram[68][55]+sumram[68][56]+sumram[68][57]+sumram[68][58]+sumram[68][59]+sumram[68][60]+sumram[68][61]+sumram[68][62]+sumram[68][63]+sumram[68][64]+sumram[68][65]+sumram[68][66]+sumram[68][67]+sumram[68][68]+sumram[68][69]+sumram[68][70]+sumram[68][71]+sumram[68][72]+sumram[68][73]+sumram[68][74]+sumram[68][75]+sumram[68][76]+sumram[68][77]+sumram[68][78]+sumram[68][79]+sumram[68][80]+sumram[68][81]+sumram[68][82]+sumram[68][83]+sumram[68][84]+sumram[68][85]+sumram[68][86]+sumram[68][87]+sumram[68][88]+sumram[68][89]+sumram[68][90]+sumram[68][91]+sumram[68][92]+sumram[68][93]+sumram[68][94]+sumram[68][95]+sumram[68][96]+sumram[68][97]+sumram[68][98]+sumram[68][99]+sumram[68][100]+sumram[68][101]+sumram[68][102]+sumram[68][103]+sumram[68][104]+sumram[68][105]+sumram[68][106]+sumram[68][107]+sumram[68][108]+sumram[68][109]+sumram[68][110]+sumram[68][111]+sumram[68][112]+sumram[68][113]+sumram[68][114]+sumram[68][115]+sumram[68][116]+sumram[68][117]+sumram[68][118]+sumram[68][119]+sumram[68][120]+sumram[68][121]+sumram[68][122]+sumram[68][123]+sumram[68][124]+sumram[68][125]+sumram[68][126]+sumram[68][127]+sumram[68][128]+sumram[68][129]+sumram[68][130]+sumram[68][131]+sumram[68][132]+sumram[68][133]+sumram[68][134]+sumram[68][135]+sumram[68][136];
    assign sumcache[69]=sumram[69][0]+sumram[69][1]+sumram[69][2]+sumram[69][3]+sumram[69][4]+sumram[69][5]+sumram[69][6]+sumram[69][7]+sumram[69][8]+sumram[69][9]+sumram[69][10]+sumram[69][11]+sumram[69][12]+sumram[69][13]+sumram[69][14]+sumram[69][15]+sumram[69][16]+sumram[69][17]+sumram[69][18]+sumram[69][19]+sumram[69][20]+sumram[69][21]+sumram[69][22]+sumram[69][23]+sumram[69][24]+sumram[69][25]+sumram[69][26]+sumram[69][27]+sumram[69][28]+sumram[69][29]+sumram[69][30]+sumram[69][31]+sumram[69][32]+sumram[69][33]+sumram[69][34]+sumram[69][35]+sumram[69][36]+sumram[69][37]+sumram[69][38]+sumram[69][39]+sumram[69][40]+sumram[69][41]+sumram[69][42]+sumram[69][43]+sumram[69][44]+sumram[69][45]+sumram[69][46]+sumram[69][47]+sumram[69][48]+sumram[69][49]+sumram[69][50]+sumram[69][51]+sumram[69][52]+sumram[69][53]+sumram[69][54]+sumram[69][55]+sumram[69][56]+sumram[69][57]+sumram[69][58]+sumram[69][59]+sumram[69][60]+sumram[69][61]+sumram[69][62]+sumram[69][63]+sumram[69][64]+sumram[69][65]+sumram[69][66]+sumram[69][67]+sumram[69][68]+sumram[69][69]+sumram[69][70]+sumram[69][71]+sumram[69][72]+sumram[69][73]+sumram[69][74]+sumram[69][75]+sumram[69][76]+sumram[69][77]+sumram[69][78]+sumram[69][79]+sumram[69][80]+sumram[69][81]+sumram[69][82]+sumram[69][83]+sumram[69][84]+sumram[69][85]+sumram[69][86]+sumram[69][87]+sumram[69][88]+sumram[69][89]+sumram[69][90]+sumram[69][91]+sumram[69][92]+sumram[69][93]+sumram[69][94]+sumram[69][95]+sumram[69][96]+sumram[69][97]+sumram[69][98]+sumram[69][99]+sumram[69][100]+sumram[69][101]+sumram[69][102]+sumram[69][103]+sumram[69][104]+sumram[69][105]+sumram[69][106]+sumram[69][107]+sumram[69][108]+sumram[69][109]+sumram[69][110]+sumram[69][111]+sumram[69][112]+sumram[69][113]+sumram[69][114]+sumram[69][115]+sumram[69][116]+sumram[69][117]+sumram[69][118]+sumram[69][119]+sumram[69][120]+sumram[69][121]+sumram[69][122]+sumram[69][123]+sumram[69][124]+sumram[69][125]+sumram[69][126]+sumram[69][127]+sumram[69][128]+sumram[69][129]+sumram[69][130]+sumram[69][131]+sumram[69][132]+sumram[69][133]+sumram[69][134]+sumram[69][135]+sumram[69][136];
    assign sumcache[70]=sumram[70][0]+sumram[70][1]+sumram[70][2]+sumram[70][3]+sumram[70][4]+sumram[70][5]+sumram[70][6]+sumram[70][7]+sumram[70][8]+sumram[70][9]+sumram[70][10]+sumram[70][11]+sumram[70][12]+sumram[70][13]+sumram[70][14]+sumram[70][15]+sumram[70][16]+sumram[70][17]+sumram[70][18]+sumram[70][19]+sumram[70][20]+sumram[70][21]+sumram[70][22]+sumram[70][23]+sumram[70][24]+sumram[70][25]+sumram[70][26]+sumram[70][27]+sumram[70][28]+sumram[70][29]+sumram[70][30]+sumram[70][31]+sumram[70][32]+sumram[70][33]+sumram[70][34]+sumram[70][35]+sumram[70][36]+sumram[70][37]+sumram[70][38]+sumram[70][39]+sumram[70][40]+sumram[70][41]+sumram[70][42]+sumram[70][43]+sumram[70][44]+sumram[70][45]+sumram[70][46]+sumram[70][47]+sumram[70][48]+sumram[70][49]+sumram[70][50]+sumram[70][51]+sumram[70][52]+sumram[70][53]+sumram[70][54]+sumram[70][55]+sumram[70][56]+sumram[70][57]+sumram[70][58]+sumram[70][59]+sumram[70][60]+sumram[70][61]+sumram[70][62]+sumram[70][63]+sumram[70][64]+sumram[70][65]+sumram[70][66]+sumram[70][67]+sumram[70][68]+sumram[70][69]+sumram[70][70]+sumram[70][71]+sumram[70][72]+sumram[70][73]+sumram[70][74]+sumram[70][75]+sumram[70][76]+sumram[70][77]+sumram[70][78]+sumram[70][79]+sumram[70][80]+sumram[70][81]+sumram[70][82]+sumram[70][83]+sumram[70][84]+sumram[70][85]+sumram[70][86]+sumram[70][87]+sumram[70][88]+sumram[70][89]+sumram[70][90]+sumram[70][91]+sumram[70][92]+sumram[70][93]+sumram[70][94]+sumram[70][95]+sumram[70][96]+sumram[70][97]+sumram[70][98]+sumram[70][99]+sumram[70][100]+sumram[70][101]+sumram[70][102]+sumram[70][103]+sumram[70][104]+sumram[70][105]+sumram[70][106]+sumram[70][107]+sumram[70][108]+sumram[70][109]+sumram[70][110]+sumram[70][111]+sumram[70][112]+sumram[70][113]+sumram[70][114]+sumram[70][115]+sumram[70][116]+sumram[70][117]+sumram[70][118]+sumram[70][119]+sumram[70][120]+sumram[70][121]+sumram[70][122]+sumram[70][123]+sumram[70][124]+sumram[70][125]+sumram[70][126]+sumram[70][127]+sumram[70][128]+sumram[70][129]+sumram[70][130]+sumram[70][131]+sumram[70][132]+sumram[70][133]+sumram[70][134]+sumram[70][135]+sumram[70][136];
    assign sumcache[71]=sumram[71][0]+sumram[71][1]+sumram[71][2]+sumram[71][3]+sumram[71][4]+sumram[71][5]+sumram[71][6]+sumram[71][7]+sumram[71][8]+sumram[71][9]+sumram[71][10]+sumram[71][11]+sumram[71][12]+sumram[71][13]+sumram[71][14]+sumram[71][15]+sumram[71][16]+sumram[71][17]+sumram[71][18]+sumram[71][19]+sumram[71][20]+sumram[71][21]+sumram[71][22]+sumram[71][23]+sumram[71][24]+sumram[71][25]+sumram[71][26]+sumram[71][27]+sumram[71][28]+sumram[71][29]+sumram[71][30]+sumram[71][31]+sumram[71][32]+sumram[71][33]+sumram[71][34]+sumram[71][35]+sumram[71][36]+sumram[71][37]+sumram[71][38]+sumram[71][39]+sumram[71][40]+sumram[71][41]+sumram[71][42]+sumram[71][43]+sumram[71][44]+sumram[71][45]+sumram[71][46]+sumram[71][47]+sumram[71][48]+sumram[71][49]+sumram[71][50]+sumram[71][51]+sumram[71][52]+sumram[71][53]+sumram[71][54]+sumram[71][55]+sumram[71][56]+sumram[71][57]+sumram[71][58]+sumram[71][59]+sumram[71][60]+sumram[71][61]+sumram[71][62]+sumram[71][63]+sumram[71][64]+sumram[71][65]+sumram[71][66]+sumram[71][67]+sumram[71][68]+sumram[71][69]+sumram[71][70]+sumram[71][71]+sumram[71][72]+sumram[71][73]+sumram[71][74]+sumram[71][75]+sumram[71][76]+sumram[71][77]+sumram[71][78]+sumram[71][79]+sumram[71][80]+sumram[71][81]+sumram[71][82]+sumram[71][83]+sumram[71][84]+sumram[71][85]+sumram[71][86]+sumram[71][87]+sumram[71][88]+sumram[71][89]+sumram[71][90]+sumram[71][91]+sumram[71][92]+sumram[71][93]+sumram[71][94]+sumram[71][95]+sumram[71][96]+sumram[71][97]+sumram[71][98]+sumram[71][99]+sumram[71][100]+sumram[71][101]+sumram[71][102]+sumram[71][103]+sumram[71][104]+sumram[71][105]+sumram[71][106]+sumram[71][107]+sumram[71][108]+sumram[71][109]+sumram[71][110]+sumram[71][111]+sumram[71][112]+sumram[71][113]+sumram[71][114]+sumram[71][115]+sumram[71][116]+sumram[71][117]+sumram[71][118]+sumram[71][119]+sumram[71][120]+sumram[71][121]+sumram[71][122]+sumram[71][123]+sumram[71][124]+sumram[71][125]+sumram[71][126]+sumram[71][127]+sumram[71][128]+sumram[71][129]+sumram[71][130]+sumram[71][131]+sumram[71][132]+sumram[71][133]+sumram[71][134]+sumram[71][135]+sumram[71][136];
    assign sumcache[72]=sumram[72][0]+sumram[72][1]+sumram[72][2]+sumram[72][3]+sumram[72][4]+sumram[72][5]+sumram[72][6]+sumram[72][7]+sumram[72][8]+sumram[72][9]+sumram[72][10]+sumram[72][11]+sumram[72][12]+sumram[72][13]+sumram[72][14]+sumram[72][15]+sumram[72][16]+sumram[72][17]+sumram[72][18]+sumram[72][19]+sumram[72][20]+sumram[72][21]+sumram[72][22]+sumram[72][23]+sumram[72][24]+sumram[72][25]+sumram[72][26]+sumram[72][27]+sumram[72][28]+sumram[72][29]+sumram[72][30]+sumram[72][31]+sumram[72][32]+sumram[72][33]+sumram[72][34]+sumram[72][35]+sumram[72][36]+sumram[72][37]+sumram[72][38]+sumram[72][39]+sumram[72][40]+sumram[72][41]+sumram[72][42]+sumram[72][43]+sumram[72][44]+sumram[72][45]+sumram[72][46]+sumram[72][47]+sumram[72][48]+sumram[72][49]+sumram[72][50]+sumram[72][51]+sumram[72][52]+sumram[72][53]+sumram[72][54]+sumram[72][55]+sumram[72][56]+sumram[72][57]+sumram[72][58]+sumram[72][59]+sumram[72][60]+sumram[72][61]+sumram[72][62]+sumram[72][63]+sumram[72][64]+sumram[72][65]+sumram[72][66]+sumram[72][67]+sumram[72][68]+sumram[72][69]+sumram[72][70]+sumram[72][71]+sumram[72][72]+sumram[72][73]+sumram[72][74]+sumram[72][75]+sumram[72][76]+sumram[72][77]+sumram[72][78]+sumram[72][79]+sumram[72][80]+sumram[72][81]+sumram[72][82]+sumram[72][83]+sumram[72][84]+sumram[72][85]+sumram[72][86]+sumram[72][87]+sumram[72][88]+sumram[72][89]+sumram[72][90]+sumram[72][91]+sumram[72][92]+sumram[72][93]+sumram[72][94]+sumram[72][95]+sumram[72][96]+sumram[72][97]+sumram[72][98]+sumram[72][99]+sumram[72][100]+sumram[72][101]+sumram[72][102]+sumram[72][103]+sumram[72][104]+sumram[72][105]+sumram[72][106]+sumram[72][107]+sumram[72][108]+sumram[72][109]+sumram[72][110]+sumram[72][111]+sumram[72][112]+sumram[72][113]+sumram[72][114]+sumram[72][115]+sumram[72][116]+sumram[72][117]+sumram[72][118]+sumram[72][119]+sumram[72][120]+sumram[72][121]+sumram[72][122]+sumram[72][123]+sumram[72][124]+sumram[72][125]+sumram[72][126]+sumram[72][127]+sumram[72][128]+sumram[72][129]+sumram[72][130]+sumram[72][131]+sumram[72][132]+sumram[72][133]+sumram[72][134]+sumram[72][135]+sumram[72][136];
    assign sumcache[73]=sumram[73][0]+sumram[73][1]+sumram[73][2]+sumram[73][3]+sumram[73][4]+sumram[73][5]+sumram[73][6]+sumram[73][7]+sumram[73][8]+sumram[73][9]+sumram[73][10]+sumram[73][11]+sumram[73][12]+sumram[73][13]+sumram[73][14]+sumram[73][15]+sumram[73][16]+sumram[73][17]+sumram[73][18]+sumram[73][19]+sumram[73][20]+sumram[73][21]+sumram[73][22]+sumram[73][23]+sumram[73][24]+sumram[73][25]+sumram[73][26]+sumram[73][27]+sumram[73][28]+sumram[73][29]+sumram[73][30]+sumram[73][31]+sumram[73][32]+sumram[73][33]+sumram[73][34]+sumram[73][35]+sumram[73][36]+sumram[73][37]+sumram[73][38]+sumram[73][39]+sumram[73][40]+sumram[73][41]+sumram[73][42]+sumram[73][43]+sumram[73][44]+sumram[73][45]+sumram[73][46]+sumram[73][47]+sumram[73][48]+sumram[73][49]+sumram[73][50]+sumram[73][51]+sumram[73][52]+sumram[73][53]+sumram[73][54]+sumram[73][55]+sumram[73][56]+sumram[73][57]+sumram[73][58]+sumram[73][59]+sumram[73][60]+sumram[73][61]+sumram[73][62]+sumram[73][63]+sumram[73][64]+sumram[73][65]+sumram[73][66]+sumram[73][67]+sumram[73][68]+sumram[73][69]+sumram[73][70]+sumram[73][71]+sumram[73][72]+sumram[73][73]+sumram[73][74]+sumram[73][75]+sumram[73][76]+sumram[73][77]+sumram[73][78]+sumram[73][79]+sumram[73][80]+sumram[73][81]+sumram[73][82]+sumram[73][83]+sumram[73][84]+sumram[73][85]+sumram[73][86]+sumram[73][87]+sumram[73][88]+sumram[73][89]+sumram[73][90]+sumram[73][91]+sumram[73][92]+sumram[73][93]+sumram[73][94]+sumram[73][95]+sumram[73][96]+sumram[73][97]+sumram[73][98]+sumram[73][99]+sumram[73][100]+sumram[73][101]+sumram[73][102]+sumram[73][103]+sumram[73][104]+sumram[73][105]+sumram[73][106]+sumram[73][107]+sumram[73][108]+sumram[73][109]+sumram[73][110]+sumram[73][111]+sumram[73][112]+sumram[73][113]+sumram[73][114]+sumram[73][115]+sumram[73][116]+sumram[73][117]+sumram[73][118]+sumram[73][119]+sumram[73][120]+sumram[73][121]+sumram[73][122]+sumram[73][123]+sumram[73][124]+sumram[73][125]+sumram[73][126]+sumram[73][127]+sumram[73][128]+sumram[73][129]+sumram[73][130]+sumram[73][131]+sumram[73][132]+sumram[73][133]+sumram[73][134]+sumram[73][135]+sumram[73][136];
    assign sumcache[74]=sumram[74][0]+sumram[74][1]+sumram[74][2]+sumram[74][3]+sumram[74][4]+sumram[74][5]+sumram[74][6]+sumram[74][7]+sumram[74][8]+sumram[74][9]+sumram[74][10]+sumram[74][11]+sumram[74][12]+sumram[74][13]+sumram[74][14]+sumram[74][15]+sumram[74][16]+sumram[74][17]+sumram[74][18]+sumram[74][19]+sumram[74][20]+sumram[74][21]+sumram[74][22]+sumram[74][23]+sumram[74][24]+sumram[74][25]+sumram[74][26]+sumram[74][27]+sumram[74][28]+sumram[74][29]+sumram[74][30]+sumram[74][31]+sumram[74][32]+sumram[74][33]+sumram[74][34]+sumram[74][35]+sumram[74][36]+sumram[74][37]+sumram[74][38]+sumram[74][39]+sumram[74][40]+sumram[74][41]+sumram[74][42]+sumram[74][43]+sumram[74][44]+sumram[74][45]+sumram[74][46]+sumram[74][47]+sumram[74][48]+sumram[74][49]+sumram[74][50]+sumram[74][51]+sumram[74][52]+sumram[74][53]+sumram[74][54]+sumram[74][55]+sumram[74][56]+sumram[74][57]+sumram[74][58]+sumram[74][59]+sumram[74][60]+sumram[74][61]+sumram[74][62]+sumram[74][63]+sumram[74][64]+sumram[74][65]+sumram[74][66]+sumram[74][67]+sumram[74][68]+sumram[74][69]+sumram[74][70]+sumram[74][71]+sumram[74][72]+sumram[74][73]+sumram[74][74]+sumram[74][75]+sumram[74][76]+sumram[74][77]+sumram[74][78]+sumram[74][79]+sumram[74][80]+sumram[74][81]+sumram[74][82]+sumram[74][83]+sumram[74][84]+sumram[74][85]+sumram[74][86]+sumram[74][87]+sumram[74][88]+sumram[74][89]+sumram[74][90]+sumram[74][91]+sumram[74][92]+sumram[74][93]+sumram[74][94]+sumram[74][95]+sumram[74][96]+sumram[74][97]+sumram[74][98]+sumram[74][99]+sumram[74][100]+sumram[74][101]+sumram[74][102]+sumram[74][103]+sumram[74][104]+sumram[74][105]+sumram[74][106]+sumram[74][107]+sumram[74][108]+sumram[74][109]+sumram[74][110]+sumram[74][111]+sumram[74][112]+sumram[74][113]+sumram[74][114]+sumram[74][115]+sumram[74][116]+sumram[74][117]+sumram[74][118]+sumram[74][119]+sumram[74][120]+sumram[74][121]+sumram[74][122]+sumram[74][123]+sumram[74][124]+sumram[74][125]+sumram[74][126]+sumram[74][127]+sumram[74][128]+sumram[74][129]+sumram[74][130]+sumram[74][131]+sumram[74][132]+sumram[74][133]+sumram[74][134]+sumram[74][135]+sumram[74][136];
    assign sumcache[75]=sumram[75][0]+sumram[75][1]+sumram[75][2]+sumram[75][3]+sumram[75][4]+sumram[75][5]+sumram[75][6]+sumram[75][7]+sumram[75][8]+sumram[75][9]+sumram[75][10]+sumram[75][11]+sumram[75][12]+sumram[75][13]+sumram[75][14]+sumram[75][15]+sumram[75][16]+sumram[75][17]+sumram[75][18]+sumram[75][19]+sumram[75][20]+sumram[75][21]+sumram[75][22]+sumram[75][23]+sumram[75][24]+sumram[75][25]+sumram[75][26]+sumram[75][27]+sumram[75][28]+sumram[75][29]+sumram[75][30]+sumram[75][31]+sumram[75][32]+sumram[75][33]+sumram[75][34]+sumram[75][35]+sumram[75][36]+sumram[75][37]+sumram[75][38]+sumram[75][39]+sumram[75][40]+sumram[75][41]+sumram[75][42]+sumram[75][43]+sumram[75][44]+sumram[75][45]+sumram[75][46]+sumram[75][47]+sumram[75][48]+sumram[75][49]+sumram[75][50]+sumram[75][51]+sumram[75][52]+sumram[75][53]+sumram[75][54]+sumram[75][55]+sumram[75][56]+sumram[75][57]+sumram[75][58]+sumram[75][59]+sumram[75][60]+sumram[75][61]+sumram[75][62]+sumram[75][63]+sumram[75][64]+sumram[75][65]+sumram[75][66]+sumram[75][67]+sumram[75][68]+sumram[75][69]+sumram[75][70]+sumram[75][71]+sumram[75][72]+sumram[75][73]+sumram[75][74]+sumram[75][75]+sumram[75][76]+sumram[75][77]+sumram[75][78]+sumram[75][79]+sumram[75][80]+sumram[75][81]+sumram[75][82]+sumram[75][83]+sumram[75][84]+sumram[75][85]+sumram[75][86]+sumram[75][87]+sumram[75][88]+sumram[75][89]+sumram[75][90]+sumram[75][91]+sumram[75][92]+sumram[75][93]+sumram[75][94]+sumram[75][95]+sumram[75][96]+sumram[75][97]+sumram[75][98]+sumram[75][99]+sumram[75][100]+sumram[75][101]+sumram[75][102]+sumram[75][103]+sumram[75][104]+sumram[75][105]+sumram[75][106]+sumram[75][107]+sumram[75][108]+sumram[75][109]+sumram[75][110]+sumram[75][111]+sumram[75][112]+sumram[75][113]+sumram[75][114]+sumram[75][115]+sumram[75][116]+sumram[75][117]+sumram[75][118]+sumram[75][119]+sumram[75][120]+sumram[75][121]+sumram[75][122]+sumram[75][123]+sumram[75][124]+sumram[75][125]+sumram[75][126]+sumram[75][127]+sumram[75][128]+sumram[75][129]+sumram[75][130]+sumram[75][131]+sumram[75][132]+sumram[75][133]+sumram[75][134]+sumram[75][135]+sumram[75][136];
    assign sumcache[76]=sumram[76][0]+sumram[76][1]+sumram[76][2]+sumram[76][3]+sumram[76][4]+sumram[76][5]+sumram[76][6]+sumram[76][7]+sumram[76][8]+sumram[76][9]+sumram[76][10]+sumram[76][11]+sumram[76][12]+sumram[76][13]+sumram[76][14]+sumram[76][15]+sumram[76][16]+sumram[76][17]+sumram[76][18]+sumram[76][19]+sumram[76][20]+sumram[76][21]+sumram[76][22]+sumram[76][23]+sumram[76][24]+sumram[76][25]+sumram[76][26]+sumram[76][27]+sumram[76][28]+sumram[76][29]+sumram[76][30]+sumram[76][31]+sumram[76][32]+sumram[76][33]+sumram[76][34]+sumram[76][35]+sumram[76][36]+sumram[76][37]+sumram[76][38]+sumram[76][39]+sumram[76][40]+sumram[76][41]+sumram[76][42]+sumram[76][43]+sumram[76][44]+sumram[76][45]+sumram[76][46]+sumram[76][47]+sumram[76][48]+sumram[76][49]+sumram[76][50]+sumram[76][51]+sumram[76][52]+sumram[76][53]+sumram[76][54]+sumram[76][55]+sumram[76][56]+sumram[76][57]+sumram[76][58]+sumram[76][59]+sumram[76][60]+sumram[76][61]+sumram[76][62]+sumram[76][63]+sumram[76][64]+sumram[76][65]+sumram[76][66]+sumram[76][67]+sumram[76][68]+sumram[76][69]+sumram[76][70]+sumram[76][71]+sumram[76][72]+sumram[76][73]+sumram[76][74]+sumram[76][75]+sumram[76][76]+sumram[76][77]+sumram[76][78]+sumram[76][79]+sumram[76][80]+sumram[76][81]+sumram[76][82]+sumram[76][83]+sumram[76][84]+sumram[76][85]+sumram[76][86]+sumram[76][87]+sumram[76][88]+sumram[76][89]+sumram[76][90]+sumram[76][91]+sumram[76][92]+sumram[76][93]+sumram[76][94]+sumram[76][95]+sumram[76][96]+sumram[76][97]+sumram[76][98]+sumram[76][99]+sumram[76][100]+sumram[76][101]+sumram[76][102]+sumram[76][103]+sumram[76][104]+sumram[76][105]+sumram[76][106]+sumram[76][107]+sumram[76][108]+sumram[76][109]+sumram[76][110]+sumram[76][111]+sumram[76][112]+sumram[76][113]+sumram[76][114]+sumram[76][115]+sumram[76][116]+sumram[76][117]+sumram[76][118]+sumram[76][119]+sumram[76][120]+sumram[76][121]+sumram[76][122]+sumram[76][123]+sumram[76][124]+sumram[76][125]+sumram[76][126]+sumram[76][127]+sumram[76][128]+sumram[76][129]+sumram[76][130]+sumram[76][131]+sumram[76][132]+sumram[76][133]+sumram[76][134]+sumram[76][135]+sumram[76][136];
    assign sumcache[77]=sumram[77][0]+sumram[77][1]+sumram[77][2]+sumram[77][3]+sumram[77][4]+sumram[77][5]+sumram[77][6]+sumram[77][7]+sumram[77][8]+sumram[77][9]+sumram[77][10]+sumram[77][11]+sumram[77][12]+sumram[77][13]+sumram[77][14]+sumram[77][15]+sumram[77][16]+sumram[77][17]+sumram[77][18]+sumram[77][19]+sumram[77][20]+sumram[77][21]+sumram[77][22]+sumram[77][23]+sumram[77][24]+sumram[77][25]+sumram[77][26]+sumram[77][27]+sumram[77][28]+sumram[77][29]+sumram[77][30]+sumram[77][31]+sumram[77][32]+sumram[77][33]+sumram[77][34]+sumram[77][35]+sumram[77][36]+sumram[77][37]+sumram[77][38]+sumram[77][39]+sumram[77][40]+sumram[77][41]+sumram[77][42]+sumram[77][43]+sumram[77][44]+sumram[77][45]+sumram[77][46]+sumram[77][47]+sumram[77][48]+sumram[77][49]+sumram[77][50]+sumram[77][51]+sumram[77][52]+sumram[77][53]+sumram[77][54]+sumram[77][55]+sumram[77][56]+sumram[77][57]+sumram[77][58]+sumram[77][59]+sumram[77][60]+sumram[77][61]+sumram[77][62]+sumram[77][63]+sumram[77][64]+sumram[77][65]+sumram[77][66]+sumram[77][67]+sumram[77][68]+sumram[77][69]+sumram[77][70]+sumram[77][71]+sumram[77][72]+sumram[77][73]+sumram[77][74]+sumram[77][75]+sumram[77][76]+sumram[77][77]+sumram[77][78]+sumram[77][79]+sumram[77][80]+sumram[77][81]+sumram[77][82]+sumram[77][83]+sumram[77][84]+sumram[77][85]+sumram[77][86]+sumram[77][87]+sumram[77][88]+sumram[77][89]+sumram[77][90]+sumram[77][91]+sumram[77][92]+sumram[77][93]+sumram[77][94]+sumram[77][95]+sumram[77][96]+sumram[77][97]+sumram[77][98]+sumram[77][99]+sumram[77][100]+sumram[77][101]+sumram[77][102]+sumram[77][103]+sumram[77][104]+sumram[77][105]+sumram[77][106]+sumram[77][107]+sumram[77][108]+sumram[77][109]+sumram[77][110]+sumram[77][111]+sumram[77][112]+sumram[77][113]+sumram[77][114]+sumram[77][115]+sumram[77][116]+sumram[77][117]+sumram[77][118]+sumram[77][119]+sumram[77][120]+sumram[77][121]+sumram[77][122]+sumram[77][123]+sumram[77][124]+sumram[77][125]+sumram[77][126]+sumram[77][127]+sumram[77][128]+sumram[77][129]+sumram[77][130]+sumram[77][131]+sumram[77][132]+sumram[77][133]+sumram[77][134]+sumram[77][135]+sumram[77][136];
    assign sumcache[78]=sumram[78][0]+sumram[78][1]+sumram[78][2]+sumram[78][3]+sumram[78][4]+sumram[78][5]+sumram[78][6]+sumram[78][7]+sumram[78][8]+sumram[78][9]+sumram[78][10]+sumram[78][11]+sumram[78][12]+sumram[78][13]+sumram[78][14]+sumram[78][15]+sumram[78][16]+sumram[78][17]+sumram[78][18]+sumram[78][19]+sumram[78][20]+sumram[78][21]+sumram[78][22]+sumram[78][23]+sumram[78][24]+sumram[78][25]+sumram[78][26]+sumram[78][27]+sumram[78][28]+sumram[78][29]+sumram[78][30]+sumram[78][31]+sumram[78][32]+sumram[78][33]+sumram[78][34]+sumram[78][35]+sumram[78][36]+sumram[78][37]+sumram[78][38]+sumram[78][39]+sumram[78][40]+sumram[78][41]+sumram[78][42]+sumram[78][43]+sumram[78][44]+sumram[78][45]+sumram[78][46]+sumram[78][47]+sumram[78][48]+sumram[78][49]+sumram[78][50]+sumram[78][51]+sumram[78][52]+sumram[78][53]+sumram[78][54]+sumram[78][55]+sumram[78][56]+sumram[78][57]+sumram[78][58]+sumram[78][59]+sumram[78][60]+sumram[78][61]+sumram[78][62]+sumram[78][63]+sumram[78][64]+sumram[78][65]+sumram[78][66]+sumram[78][67]+sumram[78][68]+sumram[78][69]+sumram[78][70]+sumram[78][71]+sumram[78][72]+sumram[78][73]+sumram[78][74]+sumram[78][75]+sumram[78][76]+sumram[78][77]+sumram[78][78]+sumram[78][79]+sumram[78][80]+sumram[78][81]+sumram[78][82]+sumram[78][83]+sumram[78][84]+sumram[78][85]+sumram[78][86]+sumram[78][87]+sumram[78][88]+sumram[78][89]+sumram[78][90]+sumram[78][91]+sumram[78][92]+sumram[78][93]+sumram[78][94]+sumram[78][95]+sumram[78][96]+sumram[78][97]+sumram[78][98]+sumram[78][99]+sumram[78][100]+sumram[78][101]+sumram[78][102]+sumram[78][103]+sumram[78][104]+sumram[78][105]+sumram[78][106]+sumram[78][107]+sumram[78][108]+sumram[78][109]+sumram[78][110]+sumram[78][111]+sumram[78][112]+sumram[78][113]+sumram[78][114]+sumram[78][115]+sumram[78][116]+sumram[78][117]+sumram[78][118]+sumram[78][119]+sumram[78][120]+sumram[78][121]+sumram[78][122]+sumram[78][123]+sumram[78][124]+sumram[78][125]+sumram[78][126]+sumram[78][127]+sumram[78][128]+sumram[78][129]+sumram[78][130]+sumram[78][131]+sumram[78][132]+sumram[78][133]+sumram[78][134]+sumram[78][135]+sumram[78][136];
    assign sumcache[79]=sumram[79][0]+sumram[79][1]+sumram[79][2]+sumram[79][3]+sumram[79][4]+sumram[79][5]+sumram[79][6]+sumram[79][7]+sumram[79][8]+sumram[79][9]+sumram[79][10]+sumram[79][11]+sumram[79][12]+sumram[79][13]+sumram[79][14]+sumram[79][15]+sumram[79][16]+sumram[79][17]+sumram[79][18]+sumram[79][19]+sumram[79][20]+sumram[79][21]+sumram[79][22]+sumram[79][23]+sumram[79][24]+sumram[79][25]+sumram[79][26]+sumram[79][27]+sumram[79][28]+sumram[79][29]+sumram[79][30]+sumram[79][31]+sumram[79][32]+sumram[79][33]+sumram[79][34]+sumram[79][35]+sumram[79][36]+sumram[79][37]+sumram[79][38]+sumram[79][39]+sumram[79][40]+sumram[79][41]+sumram[79][42]+sumram[79][43]+sumram[79][44]+sumram[79][45]+sumram[79][46]+sumram[79][47]+sumram[79][48]+sumram[79][49]+sumram[79][50]+sumram[79][51]+sumram[79][52]+sumram[79][53]+sumram[79][54]+sumram[79][55]+sumram[79][56]+sumram[79][57]+sumram[79][58]+sumram[79][59]+sumram[79][60]+sumram[79][61]+sumram[79][62]+sumram[79][63]+sumram[79][64]+sumram[79][65]+sumram[79][66]+sumram[79][67]+sumram[79][68]+sumram[79][69]+sumram[79][70]+sumram[79][71]+sumram[79][72]+sumram[79][73]+sumram[79][74]+sumram[79][75]+sumram[79][76]+sumram[79][77]+sumram[79][78]+sumram[79][79]+sumram[79][80]+sumram[79][81]+sumram[79][82]+sumram[79][83]+sumram[79][84]+sumram[79][85]+sumram[79][86]+sumram[79][87]+sumram[79][88]+sumram[79][89]+sumram[79][90]+sumram[79][91]+sumram[79][92]+sumram[79][93]+sumram[79][94]+sumram[79][95]+sumram[79][96]+sumram[79][97]+sumram[79][98]+sumram[79][99]+sumram[79][100]+sumram[79][101]+sumram[79][102]+sumram[79][103]+sumram[79][104]+sumram[79][105]+sumram[79][106]+sumram[79][107]+sumram[79][108]+sumram[79][109]+sumram[79][110]+sumram[79][111]+sumram[79][112]+sumram[79][113]+sumram[79][114]+sumram[79][115]+sumram[79][116]+sumram[79][117]+sumram[79][118]+sumram[79][119]+sumram[79][120]+sumram[79][121]+sumram[79][122]+sumram[79][123]+sumram[79][124]+sumram[79][125]+sumram[79][126]+sumram[79][127]+sumram[79][128]+sumram[79][129]+sumram[79][130]+sumram[79][131]+sumram[79][132]+sumram[79][133]+sumram[79][134]+sumram[79][135]+sumram[79][136];
    assign sumcache[80]=sumram[80][0]+sumram[80][1]+sumram[80][2]+sumram[80][3]+sumram[80][4]+sumram[80][5]+sumram[80][6]+sumram[80][7]+sumram[80][8]+sumram[80][9]+sumram[80][10]+sumram[80][11]+sumram[80][12]+sumram[80][13]+sumram[80][14]+sumram[80][15]+sumram[80][16]+sumram[80][17]+sumram[80][18]+sumram[80][19]+sumram[80][20]+sumram[80][21]+sumram[80][22]+sumram[80][23]+sumram[80][24]+sumram[80][25]+sumram[80][26]+sumram[80][27]+sumram[80][28]+sumram[80][29]+sumram[80][30]+sumram[80][31]+sumram[80][32]+sumram[80][33]+sumram[80][34]+sumram[80][35]+sumram[80][36]+sumram[80][37]+sumram[80][38]+sumram[80][39]+sumram[80][40]+sumram[80][41]+sumram[80][42]+sumram[80][43]+sumram[80][44]+sumram[80][45]+sumram[80][46]+sumram[80][47]+sumram[80][48]+sumram[80][49]+sumram[80][50]+sumram[80][51]+sumram[80][52]+sumram[80][53]+sumram[80][54]+sumram[80][55]+sumram[80][56]+sumram[80][57]+sumram[80][58]+sumram[80][59]+sumram[80][60]+sumram[80][61]+sumram[80][62]+sumram[80][63]+sumram[80][64]+sumram[80][65]+sumram[80][66]+sumram[80][67]+sumram[80][68]+sumram[80][69]+sumram[80][70]+sumram[80][71]+sumram[80][72]+sumram[80][73]+sumram[80][74]+sumram[80][75]+sumram[80][76]+sumram[80][77]+sumram[80][78]+sumram[80][79]+sumram[80][80]+sumram[80][81]+sumram[80][82]+sumram[80][83]+sumram[80][84]+sumram[80][85]+sumram[80][86]+sumram[80][87]+sumram[80][88]+sumram[80][89]+sumram[80][90]+sumram[80][91]+sumram[80][92]+sumram[80][93]+sumram[80][94]+sumram[80][95]+sumram[80][96]+sumram[80][97]+sumram[80][98]+sumram[80][99]+sumram[80][100]+sumram[80][101]+sumram[80][102]+sumram[80][103]+sumram[80][104]+sumram[80][105]+sumram[80][106]+sumram[80][107]+sumram[80][108]+sumram[80][109]+sumram[80][110]+sumram[80][111]+sumram[80][112]+sumram[80][113]+sumram[80][114]+sumram[80][115]+sumram[80][116]+sumram[80][117]+sumram[80][118]+sumram[80][119]+sumram[80][120]+sumram[80][121]+sumram[80][122]+sumram[80][123]+sumram[80][124]+sumram[80][125]+sumram[80][126]+sumram[80][127]+sumram[80][128]+sumram[80][129]+sumram[80][130]+sumram[80][131]+sumram[80][132]+sumram[80][133]+sumram[80][134]+sumram[80][135]+sumram[80][136];
    assign sumcache[81]=sumram[81][0]+sumram[81][1]+sumram[81][2]+sumram[81][3]+sumram[81][4]+sumram[81][5]+sumram[81][6]+sumram[81][7]+sumram[81][8]+sumram[81][9]+sumram[81][10]+sumram[81][11]+sumram[81][12]+sumram[81][13]+sumram[81][14]+sumram[81][15]+sumram[81][16]+sumram[81][17]+sumram[81][18]+sumram[81][19]+sumram[81][20]+sumram[81][21]+sumram[81][22]+sumram[81][23]+sumram[81][24]+sumram[81][25]+sumram[81][26]+sumram[81][27]+sumram[81][28]+sumram[81][29]+sumram[81][30]+sumram[81][31]+sumram[81][32]+sumram[81][33]+sumram[81][34]+sumram[81][35]+sumram[81][36]+sumram[81][37]+sumram[81][38]+sumram[81][39]+sumram[81][40]+sumram[81][41]+sumram[81][42]+sumram[81][43]+sumram[81][44]+sumram[81][45]+sumram[81][46]+sumram[81][47]+sumram[81][48]+sumram[81][49]+sumram[81][50]+sumram[81][51]+sumram[81][52]+sumram[81][53]+sumram[81][54]+sumram[81][55]+sumram[81][56]+sumram[81][57]+sumram[81][58]+sumram[81][59]+sumram[81][60]+sumram[81][61]+sumram[81][62]+sumram[81][63]+sumram[81][64]+sumram[81][65]+sumram[81][66]+sumram[81][67]+sumram[81][68]+sumram[81][69]+sumram[81][70]+sumram[81][71]+sumram[81][72]+sumram[81][73]+sumram[81][74]+sumram[81][75]+sumram[81][76]+sumram[81][77]+sumram[81][78]+sumram[81][79]+sumram[81][80]+sumram[81][81]+sumram[81][82]+sumram[81][83]+sumram[81][84]+sumram[81][85]+sumram[81][86]+sumram[81][87]+sumram[81][88]+sumram[81][89]+sumram[81][90]+sumram[81][91]+sumram[81][92]+sumram[81][93]+sumram[81][94]+sumram[81][95]+sumram[81][96]+sumram[81][97]+sumram[81][98]+sumram[81][99]+sumram[81][100]+sumram[81][101]+sumram[81][102]+sumram[81][103]+sumram[81][104]+sumram[81][105]+sumram[81][106]+sumram[81][107]+sumram[81][108]+sumram[81][109]+sumram[81][110]+sumram[81][111]+sumram[81][112]+sumram[81][113]+sumram[81][114]+sumram[81][115]+sumram[81][116]+sumram[81][117]+sumram[81][118]+sumram[81][119]+sumram[81][120]+sumram[81][121]+sumram[81][122]+sumram[81][123]+sumram[81][124]+sumram[81][125]+sumram[81][126]+sumram[81][127]+sumram[81][128]+sumram[81][129]+sumram[81][130]+sumram[81][131]+sumram[81][132]+sumram[81][133]+sumram[81][134]+sumram[81][135]+sumram[81][136];
    assign sumcache[82]=sumram[82][0]+sumram[82][1]+sumram[82][2]+sumram[82][3]+sumram[82][4]+sumram[82][5]+sumram[82][6]+sumram[82][7]+sumram[82][8]+sumram[82][9]+sumram[82][10]+sumram[82][11]+sumram[82][12]+sumram[82][13]+sumram[82][14]+sumram[82][15]+sumram[82][16]+sumram[82][17]+sumram[82][18]+sumram[82][19]+sumram[82][20]+sumram[82][21]+sumram[82][22]+sumram[82][23]+sumram[82][24]+sumram[82][25]+sumram[82][26]+sumram[82][27]+sumram[82][28]+sumram[82][29]+sumram[82][30]+sumram[82][31]+sumram[82][32]+sumram[82][33]+sumram[82][34]+sumram[82][35]+sumram[82][36]+sumram[82][37]+sumram[82][38]+sumram[82][39]+sumram[82][40]+sumram[82][41]+sumram[82][42]+sumram[82][43]+sumram[82][44]+sumram[82][45]+sumram[82][46]+sumram[82][47]+sumram[82][48]+sumram[82][49]+sumram[82][50]+sumram[82][51]+sumram[82][52]+sumram[82][53]+sumram[82][54]+sumram[82][55]+sumram[82][56]+sumram[82][57]+sumram[82][58]+sumram[82][59]+sumram[82][60]+sumram[82][61]+sumram[82][62]+sumram[82][63]+sumram[82][64]+sumram[82][65]+sumram[82][66]+sumram[82][67]+sumram[82][68]+sumram[82][69]+sumram[82][70]+sumram[82][71]+sumram[82][72]+sumram[82][73]+sumram[82][74]+sumram[82][75]+sumram[82][76]+sumram[82][77]+sumram[82][78]+sumram[82][79]+sumram[82][80]+sumram[82][81]+sumram[82][82]+sumram[82][83]+sumram[82][84]+sumram[82][85]+sumram[82][86]+sumram[82][87]+sumram[82][88]+sumram[82][89]+sumram[82][90]+sumram[82][91]+sumram[82][92]+sumram[82][93]+sumram[82][94]+sumram[82][95]+sumram[82][96]+sumram[82][97]+sumram[82][98]+sumram[82][99]+sumram[82][100]+sumram[82][101]+sumram[82][102]+sumram[82][103]+sumram[82][104]+sumram[82][105]+sumram[82][106]+sumram[82][107]+sumram[82][108]+sumram[82][109]+sumram[82][110]+sumram[82][111]+sumram[82][112]+sumram[82][113]+sumram[82][114]+sumram[82][115]+sumram[82][116]+sumram[82][117]+sumram[82][118]+sumram[82][119]+sumram[82][120]+sumram[82][121]+sumram[82][122]+sumram[82][123]+sumram[82][124]+sumram[82][125]+sumram[82][126]+sumram[82][127]+sumram[82][128]+sumram[82][129]+sumram[82][130]+sumram[82][131]+sumram[82][132]+sumram[82][133]+sumram[82][134]+sumram[82][135]+sumram[82][136];
    assign sumcache[83]=sumram[83][0]+sumram[83][1]+sumram[83][2]+sumram[83][3]+sumram[83][4]+sumram[83][5]+sumram[83][6]+sumram[83][7]+sumram[83][8]+sumram[83][9]+sumram[83][10]+sumram[83][11]+sumram[83][12]+sumram[83][13]+sumram[83][14]+sumram[83][15]+sumram[83][16]+sumram[83][17]+sumram[83][18]+sumram[83][19]+sumram[83][20]+sumram[83][21]+sumram[83][22]+sumram[83][23]+sumram[83][24]+sumram[83][25]+sumram[83][26]+sumram[83][27]+sumram[83][28]+sumram[83][29]+sumram[83][30]+sumram[83][31]+sumram[83][32]+sumram[83][33]+sumram[83][34]+sumram[83][35]+sumram[83][36]+sumram[83][37]+sumram[83][38]+sumram[83][39]+sumram[83][40]+sumram[83][41]+sumram[83][42]+sumram[83][43]+sumram[83][44]+sumram[83][45]+sumram[83][46]+sumram[83][47]+sumram[83][48]+sumram[83][49]+sumram[83][50]+sumram[83][51]+sumram[83][52]+sumram[83][53]+sumram[83][54]+sumram[83][55]+sumram[83][56]+sumram[83][57]+sumram[83][58]+sumram[83][59]+sumram[83][60]+sumram[83][61]+sumram[83][62]+sumram[83][63]+sumram[83][64]+sumram[83][65]+sumram[83][66]+sumram[83][67]+sumram[83][68]+sumram[83][69]+sumram[83][70]+sumram[83][71]+sumram[83][72]+sumram[83][73]+sumram[83][74]+sumram[83][75]+sumram[83][76]+sumram[83][77]+sumram[83][78]+sumram[83][79]+sumram[83][80]+sumram[83][81]+sumram[83][82]+sumram[83][83]+sumram[83][84]+sumram[83][85]+sumram[83][86]+sumram[83][87]+sumram[83][88]+sumram[83][89]+sumram[83][90]+sumram[83][91]+sumram[83][92]+sumram[83][93]+sumram[83][94]+sumram[83][95]+sumram[83][96]+sumram[83][97]+sumram[83][98]+sumram[83][99]+sumram[83][100]+sumram[83][101]+sumram[83][102]+sumram[83][103]+sumram[83][104]+sumram[83][105]+sumram[83][106]+sumram[83][107]+sumram[83][108]+sumram[83][109]+sumram[83][110]+sumram[83][111]+sumram[83][112]+sumram[83][113]+sumram[83][114]+sumram[83][115]+sumram[83][116]+sumram[83][117]+sumram[83][118]+sumram[83][119]+sumram[83][120]+sumram[83][121]+sumram[83][122]+sumram[83][123]+sumram[83][124]+sumram[83][125]+sumram[83][126]+sumram[83][127]+sumram[83][128]+sumram[83][129]+sumram[83][130]+sumram[83][131]+sumram[83][132]+sumram[83][133]+sumram[83][134]+sumram[83][135]+sumram[83][136];
    assign sumcache[84]=sumram[84][0]+sumram[84][1]+sumram[84][2]+sumram[84][3]+sumram[84][4]+sumram[84][5]+sumram[84][6]+sumram[84][7]+sumram[84][8]+sumram[84][9]+sumram[84][10]+sumram[84][11]+sumram[84][12]+sumram[84][13]+sumram[84][14]+sumram[84][15]+sumram[84][16]+sumram[84][17]+sumram[84][18]+sumram[84][19]+sumram[84][20]+sumram[84][21]+sumram[84][22]+sumram[84][23]+sumram[84][24]+sumram[84][25]+sumram[84][26]+sumram[84][27]+sumram[84][28]+sumram[84][29]+sumram[84][30]+sumram[84][31]+sumram[84][32]+sumram[84][33]+sumram[84][34]+sumram[84][35]+sumram[84][36]+sumram[84][37]+sumram[84][38]+sumram[84][39]+sumram[84][40]+sumram[84][41]+sumram[84][42]+sumram[84][43]+sumram[84][44]+sumram[84][45]+sumram[84][46]+sumram[84][47]+sumram[84][48]+sumram[84][49]+sumram[84][50]+sumram[84][51]+sumram[84][52]+sumram[84][53]+sumram[84][54]+sumram[84][55]+sumram[84][56]+sumram[84][57]+sumram[84][58]+sumram[84][59]+sumram[84][60]+sumram[84][61]+sumram[84][62]+sumram[84][63]+sumram[84][64]+sumram[84][65]+sumram[84][66]+sumram[84][67]+sumram[84][68]+sumram[84][69]+sumram[84][70]+sumram[84][71]+sumram[84][72]+sumram[84][73]+sumram[84][74]+sumram[84][75]+sumram[84][76]+sumram[84][77]+sumram[84][78]+sumram[84][79]+sumram[84][80]+sumram[84][81]+sumram[84][82]+sumram[84][83]+sumram[84][84]+sumram[84][85]+sumram[84][86]+sumram[84][87]+sumram[84][88]+sumram[84][89]+sumram[84][90]+sumram[84][91]+sumram[84][92]+sumram[84][93]+sumram[84][94]+sumram[84][95]+sumram[84][96]+sumram[84][97]+sumram[84][98]+sumram[84][99]+sumram[84][100]+sumram[84][101]+sumram[84][102]+sumram[84][103]+sumram[84][104]+sumram[84][105]+sumram[84][106]+sumram[84][107]+sumram[84][108]+sumram[84][109]+sumram[84][110]+sumram[84][111]+sumram[84][112]+sumram[84][113]+sumram[84][114]+sumram[84][115]+sumram[84][116]+sumram[84][117]+sumram[84][118]+sumram[84][119]+sumram[84][120]+sumram[84][121]+sumram[84][122]+sumram[84][123]+sumram[84][124]+sumram[84][125]+sumram[84][126]+sumram[84][127]+sumram[84][128]+sumram[84][129]+sumram[84][130]+sumram[84][131]+sumram[84][132]+sumram[84][133]+sumram[84][134]+sumram[84][135]+sumram[84][136];
    assign sumcache[85]=sumram[85][0]+sumram[85][1]+sumram[85][2]+sumram[85][3]+sumram[85][4]+sumram[85][5]+sumram[85][6]+sumram[85][7]+sumram[85][8]+sumram[85][9]+sumram[85][10]+sumram[85][11]+sumram[85][12]+sumram[85][13]+sumram[85][14]+sumram[85][15]+sumram[85][16]+sumram[85][17]+sumram[85][18]+sumram[85][19]+sumram[85][20]+sumram[85][21]+sumram[85][22]+sumram[85][23]+sumram[85][24]+sumram[85][25]+sumram[85][26]+sumram[85][27]+sumram[85][28]+sumram[85][29]+sumram[85][30]+sumram[85][31]+sumram[85][32]+sumram[85][33]+sumram[85][34]+sumram[85][35]+sumram[85][36]+sumram[85][37]+sumram[85][38]+sumram[85][39]+sumram[85][40]+sumram[85][41]+sumram[85][42]+sumram[85][43]+sumram[85][44]+sumram[85][45]+sumram[85][46]+sumram[85][47]+sumram[85][48]+sumram[85][49]+sumram[85][50]+sumram[85][51]+sumram[85][52]+sumram[85][53]+sumram[85][54]+sumram[85][55]+sumram[85][56]+sumram[85][57]+sumram[85][58]+sumram[85][59]+sumram[85][60]+sumram[85][61]+sumram[85][62]+sumram[85][63]+sumram[85][64]+sumram[85][65]+sumram[85][66]+sumram[85][67]+sumram[85][68]+sumram[85][69]+sumram[85][70]+sumram[85][71]+sumram[85][72]+sumram[85][73]+sumram[85][74]+sumram[85][75]+sumram[85][76]+sumram[85][77]+sumram[85][78]+sumram[85][79]+sumram[85][80]+sumram[85][81]+sumram[85][82]+sumram[85][83]+sumram[85][84]+sumram[85][85]+sumram[85][86]+sumram[85][87]+sumram[85][88]+sumram[85][89]+sumram[85][90]+sumram[85][91]+sumram[85][92]+sumram[85][93]+sumram[85][94]+sumram[85][95]+sumram[85][96]+sumram[85][97]+sumram[85][98]+sumram[85][99]+sumram[85][100]+sumram[85][101]+sumram[85][102]+sumram[85][103]+sumram[85][104]+sumram[85][105]+sumram[85][106]+sumram[85][107]+sumram[85][108]+sumram[85][109]+sumram[85][110]+sumram[85][111]+sumram[85][112]+sumram[85][113]+sumram[85][114]+sumram[85][115]+sumram[85][116]+sumram[85][117]+sumram[85][118]+sumram[85][119]+sumram[85][120]+sumram[85][121]+sumram[85][122]+sumram[85][123]+sumram[85][124]+sumram[85][125]+sumram[85][126]+sumram[85][127]+sumram[85][128]+sumram[85][129]+sumram[85][130]+sumram[85][131]+sumram[85][132]+sumram[85][133]+sumram[85][134]+sumram[85][135]+sumram[85][136];
    assign sumcache[86]=sumram[86][0]+sumram[86][1]+sumram[86][2]+sumram[86][3]+sumram[86][4]+sumram[86][5]+sumram[86][6]+sumram[86][7]+sumram[86][8]+sumram[86][9]+sumram[86][10]+sumram[86][11]+sumram[86][12]+sumram[86][13]+sumram[86][14]+sumram[86][15]+sumram[86][16]+sumram[86][17]+sumram[86][18]+sumram[86][19]+sumram[86][20]+sumram[86][21]+sumram[86][22]+sumram[86][23]+sumram[86][24]+sumram[86][25]+sumram[86][26]+sumram[86][27]+sumram[86][28]+sumram[86][29]+sumram[86][30]+sumram[86][31]+sumram[86][32]+sumram[86][33]+sumram[86][34]+sumram[86][35]+sumram[86][36]+sumram[86][37]+sumram[86][38]+sumram[86][39]+sumram[86][40]+sumram[86][41]+sumram[86][42]+sumram[86][43]+sumram[86][44]+sumram[86][45]+sumram[86][46]+sumram[86][47]+sumram[86][48]+sumram[86][49]+sumram[86][50]+sumram[86][51]+sumram[86][52]+sumram[86][53]+sumram[86][54]+sumram[86][55]+sumram[86][56]+sumram[86][57]+sumram[86][58]+sumram[86][59]+sumram[86][60]+sumram[86][61]+sumram[86][62]+sumram[86][63]+sumram[86][64]+sumram[86][65]+sumram[86][66]+sumram[86][67]+sumram[86][68]+sumram[86][69]+sumram[86][70]+sumram[86][71]+sumram[86][72]+sumram[86][73]+sumram[86][74]+sumram[86][75]+sumram[86][76]+sumram[86][77]+sumram[86][78]+sumram[86][79]+sumram[86][80]+sumram[86][81]+sumram[86][82]+sumram[86][83]+sumram[86][84]+sumram[86][85]+sumram[86][86]+sumram[86][87]+sumram[86][88]+sumram[86][89]+sumram[86][90]+sumram[86][91]+sumram[86][92]+sumram[86][93]+sumram[86][94]+sumram[86][95]+sumram[86][96]+sumram[86][97]+sumram[86][98]+sumram[86][99]+sumram[86][100]+sumram[86][101]+sumram[86][102]+sumram[86][103]+sumram[86][104]+sumram[86][105]+sumram[86][106]+sumram[86][107]+sumram[86][108]+sumram[86][109]+sumram[86][110]+sumram[86][111]+sumram[86][112]+sumram[86][113]+sumram[86][114]+sumram[86][115]+sumram[86][116]+sumram[86][117]+sumram[86][118]+sumram[86][119]+sumram[86][120]+sumram[86][121]+sumram[86][122]+sumram[86][123]+sumram[86][124]+sumram[86][125]+sumram[86][126]+sumram[86][127]+sumram[86][128]+sumram[86][129]+sumram[86][130]+sumram[86][131]+sumram[86][132]+sumram[86][133]+sumram[86][134]+sumram[86][135]+sumram[86][136];
    assign sumcache[87]=sumram[87][0]+sumram[87][1]+sumram[87][2]+sumram[87][3]+sumram[87][4]+sumram[87][5]+sumram[87][6]+sumram[87][7]+sumram[87][8]+sumram[87][9]+sumram[87][10]+sumram[87][11]+sumram[87][12]+sumram[87][13]+sumram[87][14]+sumram[87][15]+sumram[87][16]+sumram[87][17]+sumram[87][18]+sumram[87][19]+sumram[87][20]+sumram[87][21]+sumram[87][22]+sumram[87][23]+sumram[87][24]+sumram[87][25]+sumram[87][26]+sumram[87][27]+sumram[87][28]+sumram[87][29]+sumram[87][30]+sumram[87][31]+sumram[87][32]+sumram[87][33]+sumram[87][34]+sumram[87][35]+sumram[87][36]+sumram[87][37]+sumram[87][38]+sumram[87][39]+sumram[87][40]+sumram[87][41]+sumram[87][42]+sumram[87][43]+sumram[87][44]+sumram[87][45]+sumram[87][46]+sumram[87][47]+sumram[87][48]+sumram[87][49]+sumram[87][50]+sumram[87][51]+sumram[87][52]+sumram[87][53]+sumram[87][54]+sumram[87][55]+sumram[87][56]+sumram[87][57]+sumram[87][58]+sumram[87][59]+sumram[87][60]+sumram[87][61]+sumram[87][62]+sumram[87][63]+sumram[87][64]+sumram[87][65]+sumram[87][66]+sumram[87][67]+sumram[87][68]+sumram[87][69]+sumram[87][70]+sumram[87][71]+sumram[87][72]+sumram[87][73]+sumram[87][74]+sumram[87][75]+sumram[87][76]+sumram[87][77]+sumram[87][78]+sumram[87][79]+sumram[87][80]+sumram[87][81]+sumram[87][82]+sumram[87][83]+sumram[87][84]+sumram[87][85]+sumram[87][86]+sumram[87][87]+sumram[87][88]+sumram[87][89]+sumram[87][90]+sumram[87][91]+sumram[87][92]+sumram[87][93]+sumram[87][94]+sumram[87][95]+sumram[87][96]+sumram[87][97]+sumram[87][98]+sumram[87][99]+sumram[87][100]+sumram[87][101]+sumram[87][102]+sumram[87][103]+sumram[87][104]+sumram[87][105]+sumram[87][106]+sumram[87][107]+sumram[87][108]+sumram[87][109]+sumram[87][110]+sumram[87][111]+sumram[87][112]+sumram[87][113]+sumram[87][114]+sumram[87][115]+sumram[87][116]+sumram[87][117]+sumram[87][118]+sumram[87][119]+sumram[87][120]+sumram[87][121]+sumram[87][122]+sumram[87][123]+sumram[87][124]+sumram[87][125]+sumram[87][126]+sumram[87][127]+sumram[87][128]+sumram[87][129]+sumram[87][130]+sumram[87][131]+sumram[87][132]+sumram[87][133]+sumram[87][134]+sumram[87][135]+sumram[87][136];
    assign sumcache[88]=sumram[88][0]+sumram[88][1]+sumram[88][2]+sumram[88][3]+sumram[88][4]+sumram[88][5]+sumram[88][6]+sumram[88][7]+sumram[88][8]+sumram[88][9]+sumram[88][10]+sumram[88][11]+sumram[88][12]+sumram[88][13]+sumram[88][14]+sumram[88][15]+sumram[88][16]+sumram[88][17]+sumram[88][18]+sumram[88][19]+sumram[88][20]+sumram[88][21]+sumram[88][22]+sumram[88][23]+sumram[88][24]+sumram[88][25]+sumram[88][26]+sumram[88][27]+sumram[88][28]+sumram[88][29]+sumram[88][30]+sumram[88][31]+sumram[88][32]+sumram[88][33]+sumram[88][34]+sumram[88][35]+sumram[88][36]+sumram[88][37]+sumram[88][38]+sumram[88][39]+sumram[88][40]+sumram[88][41]+sumram[88][42]+sumram[88][43]+sumram[88][44]+sumram[88][45]+sumram[88][46]+sumram[88][47]+sumram[88][48]+sumram[88][49]+sumram[88][50]+sumram[88][51]+sumram[88][52]+sumram[88][53]+sumram[88][54]+sumram[88][55]+sumram[88][56]+sumram[88][57]+sumram[88][58]+sumram[88][59]+sumram[88][60]+sumram[88][61]+sumram[88][62]+sumram[88][63]+sumram[88][64]+sumram[88][65]+sumram[88][66]+sumram[88][67]+sumram[88][68]+sumram[88][69]+sumram[88][70]+sumram[88][71]+sumram[88][72]+sumram[88][73]+sumram[88][74]+sumram[88][75]+sumram[88][76]+sumram[88][77]+sumram[88][78]+sumram[88][79]+sumram[88][80]+sumram[88][81]+sumram[88][82]+sumram[88][83]+sumram[88][84]+sumram[88][85]+sumram[88][86]+sumram[88][87]+sumram[88][88]+sumram[88][89]+sumram[88][90]+sumram[88][91]+sumram[88][92]+sumram[88][93]+sumram[88][94]+sumram[88][95]+sumram[88][96]+sumram[88][97]+sumram[88][98]+sumram[88][99]+sumram[88][100]+sumram[88][101]+sumram[88][102]+sumram[88][103]+sumram[88][104]+sumram[88][105]+sumram[88][106]+sumram[88][107]+sumram[88][108]+sumram[88][109]+sumram[88][110]+sumram[88][111]+sumram[88][112]+sumram[88][113]+sumram[88][114]+sumram[88][115]+sumram[88][116]+sumram[88][117]+sumram[88][118]+sumram[88][119]+sumram[88][120]+sumram[88][121]+sumram[88][122]+sumram[88][123]+sumram[88][124]+sumram[88][125]+sumram[88][126]+sumram[88][127]+sumram[88][128]+sumram[88][129]+sumram[88][130]+sumram[88][131]+sumram[88][132]+sumram[88][133]+sumram[88][134]+sumram[88][135]+sumram[88][136];
    assign sumcache[89]=sumram[89][0]+sumram[89][1]+sumram[89][2]+sumram[89][3]+sumram[89][4]+sumram[89][5]+sumram[89][6]+sumram[89][7]+sumram[89][8]+sumram[89][9]+sumram[89][10]+sumram[89][11]+sumram[89][12]+sumram[89][13]+sumram[89][14]+sumram[89][15]+sumram[89][16]+sumram[89][17]+sumram[89][18]+sumram[89][19]+sumram[89][20]+sumram[89][21]+sumram[89][22]+sumram[89][23]+sumram[89][24]+sumram[89][25]+sumram[89][26]+sumram[89][27]+sumram[89][28]+sumram[89][29]+sumram[89][30]+sumram[89][31]+sumram[89][32]+sumram[89][33]+sumram[89][34]+sumram[89][35]+sumram[89][36]+sumram[89][37]+sumram[89][38]+sumram[89][39]+sumram[89][40]+sumram[89][41]+sumram[89][42]+sumram[89][43]+sumram[89][44]+sumram[89][45]+sumram[89][46]+sumram[89][47]+sumram[89][48]+sumram[89][49]+sumram[89][50]+sumram[89][51]+sumram[89][52]+sumram[89][53]+sumram[89][54]+sumram[89][55]+sumram[89][56]+sumram[89][57]+sumram[89][58]+sumram[89][59]+sumram[89][60]+sumram[89][61]+sumram[89][62]+sumram[89][63]+sumram[89][64]+sumram[89][65]+sumram[89][66]+sumram[89][67]+sumram[89][68]+sumram[89][69]+sumram[89][70]+sumram[89][71]+sumram[89][72]+sumram[89][73]+sumram[89][74]+sumram[89][75]+sumram[89][76]+sumram[89][77]+sumram[89][78]+sumram[89][79]+sumram[89][80]+sumram[89][81]+sumram[89][82]+sumram[89][83]+sumram[89][84]+sumram[89][85]+sumram[89][86]+sumram[89][87]+sumram[89][88]+sumram[89][89]+sumram[89][90]+sumram[89][91]+sumram[89][92]+sumram[89][93]+sumram[89][94]+sumram[89][95]+sumram[89][96]+sumram[89][97]+sumram[89][98]+sumram[89][99]+sumram[89][100]+sumram[89][101]+sumram[89][102]+sumram[89][103]+sumram[89][104]+sumram[89][105]+sumram[89][106]+sumram[89][107]+sumram[89][108]+sumram[89][109]+sumram[89][110]+sumram[89][111]+sumram[89][112]+sumram[89][113]+sumram[89][114]+sumram[89][115]+sumram[89][116]+sumram[89][117]+sumram[89][118]+sumram[89][119]+sumram[89][120]+sumram[89][121]+sumram[89][122]+sumram[89][123]+sumram[89][124]+sumram[89][125]+sumram[89][126]+sumram[89][127]+sumram[89][128]+sumram[89][129]+sumram[89][130]+sumram[89][131]+sumram[89][132]+sumram[89][133]+sumram[89][134]+sumram[89][135]+sumram[89][136];
    assign sumcache[90]=sumram[90][0]+sumram[90][1]+sumram[90][2]+sumram[90][3]+sumram[90][4]+sumram[90][5]+sumram[90][6]+sumram[90][7]+sumram[90][8]+sumram[90][9]+sumram[90][10]+sumram[90][11]+sumram[90][12]+sumram[90][13]+sumram[90][14]+sumram[90][15]+sumram[90][16]+sumram[90][17]+sumram[90][18]+sumram[90][19]+sumram[90][20]+sumram[90][21]+sumram[90][22]+sumram[90][23]+sumram[90][24]+sumram[90][25]+sumram[90][26]+sumram[90][27]+sumram[90][28]+sumram[90][29]+sumram[90][30]+sumram[90][31]+sumram[90][32]+sumram[90][33]+sumram[90][34]+sumram[90][35]+sumram[90][36]+sumram[90][37]+sumram[90][38]+sumram[90][39]+sumram[90][40]+sumram[90][41]+sumram[90][42]+sumram[90][43]+sumram[90][44]+sumram[90][45]+sumram[90][46]+sumram[90][47]+sumram[90][48]+sumram[90][49]+sumram[90][50]+sumram[90][51]+sumram[90][52]+sumram[90][53]+sumram[90][54]+sumram[90][55]+sumram[90][56]+sumram[90][57]+sumram[90][58]+sumram[90][59]+sumram[90][60]+sumram[90][61]+sumram[90][62]+sumram[90][63]+sumram[90][64]+sumram[90][65]+sumram[90][66]+sumram[90][67]+sumram[90][68]+sumram[90][69]+sumram[90][70]+sumram[90][71]+sumram[90][72]+sumram[90][73]+sumram[90][74]+sumram[90][75]+sumram[90][76]+sumram[90][77]+sumram[90][78]+sumram[90][79]+sumram[90][80]+sumram[90][81]+sumram[90][82]+sumram[90][83]+sumram[90][84]+sumram[90][85]+sumram[90][86]+sumram[90][87]+sumram[90][88]+sumram[90][89]+sumram[90][90]+sumram[90][91]+sumram[90][92]+sumram[90][93]+sumram[90][94]+sumram[90][95]+sumram[90][96]+sumram[90][97]+sumram[90][98]+sumram[90][99]+sumram[90][100]+sumram[90][101]+sumram[90][102]+sumram[90][103]+sumram[90][104]+sumram[90][105]+sumram[90][106]+sumram[90][107]+sumram[90][108]+sumram[90][109]+sumram[90][110]+sumram[90][111]+sumram[90][112]+sumram[90][113]+sumram[90][114]+sumram[90][115]+sumram[90][116]+sumram[90][117]+sumram[90][118]+sumram[90][119]+sumram[90][120]+sumram[90][121]+sumram[90][122]+sumram[90][123]+sumram[90][124]+sumram[90][125]+sumram[90][126]+sumram[90][127]+sumram[90][128]+sumram[90][129]+sumram[90][130]+sumram[90][131]+sumram[90][132]+sumram[90][133]+sumram[90][134]+sumram[90][135]+sumram[90][136];
    assign sumcache[91]=sumram[91][0]+sumram[91][1]+sumram[91][2]+sumram[91][3]+sumram[91][4]+sumram[91][5]+sumram[91][6]+sumram[91][7]+sumram[91][8]+sumram[91][9]+sumram[91][10]+sumram[91][11]+sumram[91][12]+sumram[91][13]+sumram[91][14]+sumram[91][15]+sumram[91][16]+sumram[91][17]+sumram[91][18]+sumram[91][19]+sumram[91][20]+sumram[91][21]+sumram[91][22]+sumram[91][23]+sumram[91][24]+sumram[91][25]+sumram[91][26]+sumram[91][27]+sumram[91][28]+sumram[91][29]+sumram[91][30]+sumram[91][31]+sumram[91][32]+sumram[91][33]+sumram[91][34]+sumram[91][35]+sumram[91][36]+sumram[91][37]+sumram[91][38]+sumram[91][39]+sumram[91][40]+sumram[91][41]+sumram[91][42]+sumram[91][43]+sumram[91][44]+sumram[91][45]+sumram[91][46]+sumram[91][47]+sumram[91][48]+sumram[91][49]+sumram[91][50]+sumram[91][51]+sumram[91][52]+sumram[91][53]+sumram[91][54]+sumram[91][55]+sumram[91][56]+sumram[91][57]+sumram[91][58]+sumram[91][59]+sumram[91][60]+sumram[91][61]+sumram[91][62]+sumram[91][63]+sumram[91][64]+sumram[91][65]+sumram[91][66]+sumram[91][67]+sumram[91][68]+sumram[91][69]+sumram[91][70]+sumram[91][71]+sumram[91][72]+sumram[91][73]+sumram[91][74]+sumram[91][75]+sumram[91][76]+sumram[91][77]+sumram[91][78]+sumram[91][79]+sumram[91][80]+sumram[91][81]+sumram[91][82]+sumram[91][83]+sumram[91][84]+sumram[91][85]+sumram[91][86]+sumram[91][87]+sumram[91][88]+sumram[91][89]+sumram[91][90]+sumram[91][91]+sumram[91][92]+sumram[91][93]+sumram[91][94]+sumram[91][95]+sumram[91][96]+sumram[91][97]+sumram[91][98]+sumram[91][99]+sumram[91][100]+sumram[91][101]+sumram[91][102]+sumram[91][103]+sumram[91][104]+sumram[91][105]+sumram[91][106]+sumram[91][107]+sumram[91][108]+sumram[91][109]+sumram[91][110]+sumram[91][111]+sumram[91][112]+sumram[91][113]+sumram[91][114]+sumram[91][115]+sumram[91][116]+sumram[91][117]+sumram[91][118]+sumram[91][119]+sumram[91][120]+sumram[91][121]+sumram[91][122]+sumram[91][123]+sumram[91][124]+sumram[91][125]+sumram[91][126]+sumram[91][127]+sumram[91][128]+sumram[91][129]+sumram[91][130]+sumram[91][131]+sumram[91][132]+sumram[91][133]+sumram[91][134]+sumram[91][135]+sumram[91][136];
    assign sumcache[92]=sumram[92][0]+sumram[92][1]+sumram[92][2]+sumram[92][3]+sumram[92][4]+sumram[92][5]+sumram[92][6]+sumram[92][7]+sumram[92][8]+sumram[92][9]+sumram[92][10]+sumram[92][11]+sumram[92][12]+sumram[92][13]+sumram[92][14]+sumram[92][15]+sumram[92][16]+sumram[92][17]+sumram[92][18]+sumram[92][19]+sumram[92][20]+sumram[92][21]+sumram[92][22]+sumram[92][23]+sumram[92][24]+sumram[92][25]+sumram[92][26]+sumram[92][27]+sumram[92][28]+sumram[92][29]+sumram[92][30]+sumram[92][31]+sumram[92][32]+sumram[92][33]+sumram[92][34]+sumram[92][35]+sumram[92][36]+sumram[92][37]+sumram[92][38]+sumram[92][39]+sumram[92][40]+sumram[92][41]+sumram[92][42]+sumram[92][43]+sumram[92][44]+sumram[92][45]+sumram[92][46]+sumram[92][47]+sumram[92][48]+sumram[92][49]+sumram[92][50]+sumram[92][51]+sumram[92][52]+sumram[92][53]+sumram[92][54]+sumram[92][55]+sumram[92][56]+sumram[92][57]+sumram[92][58]+sumram[92][59]+sumram[92][60]+sumram[92][61]+sumram[92][62]+sumram[92][63]+sumram[92][64]+sumram[92][65]+sumram[92][66]+sumram[92][67]+sumram[92][68]+sumram[92][69]+sumram[92][70]+sumram[92][71]+sumram[92][72]+sumram[92][73]+sumram[92][74]+sumram[92][75]+sumram[92][76]+sumram[92][77]+sumram[92][78]+sumram[92][79]+sumram[92][80]+sumram[92][81]+sumram[92][82]+sumram[92][83]+sumram[92][84]+sumram[92][85]+sumram[92][86]+sumram[92][87]+sumram[92][88]+sumram[92][89]+sumram[92][90]+sumram[92][91]+sumram[92][92]+sumram[92][93]+sumram[92][94]+sumram[92][95]+sumram[92][96]+sumram[92][97]+sumram[92][98]+sumram[92][99]+sumram[92][100]+sumram[92][101]+sumram[92][102]+sumram[92][103]+sumram[92][104]+sumram[92][105]+sumram[92][106]+sumram[92][107]+sumram[92][108]+sumram[92][109]+sumram[92][110]+sumram[92][111]+sumram[92][112]+sumram[92][113]+sumram[92][114]+sumram[92][115]+sumram[92][116]+sumram[92][117]+sumram[92][118]+sumram[92][119]+sumram[92][120]+sumram[92][121]+sumram[92][122]+sumram[92][123]+sumram[92][124]+sumram[92][125]+sumram[92][126]+sumram[92][127]+sumram[92][128]+sumram[92][129]+sumram[92][130]+sumram[92][131]+sumram[92][132]+sumram[92][133]+sumram[92][134]+sumram[92][135]+sumram[92][136];
    assign sumcache[93]=sumram[93][0]+sumram[93][1]+sumram[93][2]+sumram[93][3]+sumram[93][4]+sumram[93][5]+sumram[93][6]+sumram[93][7]+sumram[93][8]+sumram[93][9]+sumram[93][10]+sumram[93][11]+sumram[93][12]+sumram[93][13]+sumram[93][14]+sumram[93][15]+sumram[93][16]+sumram[93][17]+sumram[93][18]+sumram[93][19]+sumram[93][20]+sumram[93][21]+sumram[93][22]+sumram[93][23]+sumram[93][24]+sumram[93][25]+sumram[93][26]+sumram[93][27]+sumram[93][28]+sumram[93][29]+sumram[93][30]+sumram[93][31]+sumram[93][32]+sumram[93][33]+sumram[93][34]+sumram[93][35]+sumram[93][36]+sumram[93][37]+sumram[93][38]+sumram[93][39]+sumram[93][40]+sumram[93][41]+sumram[93][42]+sumram[93][43]+sumram[93][44]+sumram[93][45]+sumram[93][46]+sumram[93][47]+sumram[93][48]+sumram[93][49]+sumram[93][50]+sumram[93][51]+sumram[93][52]+sumram[93][53]+sumram[93][54]+sumram[93][55]+sumram[93][56]+sumram[93][57]+sumram[93][58]+sumram[93][59]+sumram[93][60]+sumram[93][61]+sumram[93][62]+sumram[93][63]+sumram[93][64]+sumram[93][65]+sumram[93][66]+sumram[93][67]+sumram[93][68]+sumram[93][69]+sumram[93][70]+sumram[93][71]+sumram[93][72]+sumram[93][73]+sumram[93][74]+sumram[93][75]+sumram[93][76]+sumram[93][77]+sumram[93][78]+sumram[93][79]+sumram[93][80]+sumram[93][81]+sumram[93][82]+sumram[93][83]+sumram[93][84]+sumram[93][85]+sumram[93][86]+sumram[93][87]+sumram[93][88]+sumram[93][89]+sumram[93][90]+sumram[93][91]+sumram[93][92]+sumram[93][93]+sumram[93][94]+sumram[93][95]+sumram[93][96]+sumram[93][97]+sumram[93][98]+sumram[93][99]+sumram[93][100]+sumram[93][101]+sumram[93][102]+sumram[93][103]+sumram[93][104]+sumram[93][105]+sumram[93][106]+sumram[93][107]+sumram[93][108]+sumram[93][109]+sumram[93][110]+sumram[93][111]+sumram[93][112]+sumram[93][113]+sumram[93][114]+sumram[93][115]+sumram[93][116]+sumram[93][117]+sumram[93][118]+sumram[93][119]+sumram[93][120]+sumram[93][121]+sumram[93][122]+sumram[93][123]+sumram[93][124]+sumram[93][125]+sumram[93][126]+sumram[93][127]+sumram[93][128]+sumram[93][129]+sumram[93][130]+sumram[93][131]+sumram[93][132]+sumram[93][133]+sumram[93][134]+sumram[93][135]+sumram[93][136];
    assign sumcache[94]=sumram[94][0]+sumram[94][1]+sumram[94][2]+sumram[94][3]+sumram[94][4]+sumram[94][5]+sumram[94][6]+sumram[94][7]+sumram[94][8]+sumram[94][9]+sumram[94][10]+sumram[94][11]+sumram[94][12]+sumram[94][13]+sumram[94][14]+sumram[94][15]+sumram[94][16]+sumram[94][17]+sumram[94][18]+sumram[94][19]+sumram[94][20]+sumram[94][21]+sumram[94][22]+sumram[94][23]+sumram[94][24]+sumram[94][25]+sumram[94][26]+sumram[94][27]+sumram[94][28]+sumram[94][29]+sumram[94][30]+sumram[94][31]+sumram[94][32]+sumram[94][33]+sumram[94][34]+sumram[94][35]+sumram[94][36]+sumram[94][37]+sumram[94][38]+sumram[94][39]+sumram[94][40]+sumram[94][41]+sumram[94][42]+sumram[94][43]+sumram[94][44]+sumram[94][45]+sumram[94][46]+sumram[94][47]+sumram[94][48]+sumram[94][49]+sumram[94][50]+sumram[94][51]+sumram[94][52]+sumram[94][53]+sumram[94][54]+sumram[94][55]+sumram[94][56]+sumram[94][57]+sumram[94][58]+sumram[94][59]+sumram[94][60]+sumram[94][61]+sumram[94][62]+sumram[94][63]+sumram[94][64]+sumram[94][65]+sumram[94][66]+sumram[94][67]+sumram[94][68]+sumram[94][69]+sumram[94][70]+sumram[94][71]+sumram[94][72]+sumram[94][73]+sumram[94][74]+sumram[94][75]+sumram[94][76]+sumram[94][77]+sumram[94][78]+sumram[94][79]+sumram[94][80]+sumram[94][81]+sumram[94][82]+sumram[94][83]+sumram[94][84]+sumram[94][85]+sumram[94][86]+sumram[94][87]+sumram[94][88]+sumram[94][89]+sumram[94][90]+sumram[94][91]+sumram[94][92]+sumram[94][93]+sumram[94][94]+sumram[94][95]+sumram[94][96]+sumram[94][97]+sumram[94][98]+sumram[94][99]+sumram[94][100]+sumram[94][101]+sumram[94][102]+sumram[94][103]+sumram[94][104]+sumram[94][105]+sumram[94][106]+sumram[94][107]+sumram[94][108]+sumram[94][109]+sumram[94][110]+sumram[94][111]+sumram[94][112]+sumram[94][113]+sumram[94][114]+sumram[94][115]+sumram[94][116]+sumram[94][117]+sumram[94][118]+sumram[94][119]+sumram[94][120]+sumram[94][121]+sumram[94][122]+sumram[94][123]+sumram[94][124]+sumram[94][125]+sumram[94][126]+sumram[94][127]+sumram[94][128]+sumram[94][129]+sumram[94][130]+sumram[94][131]+sumram[94][132]+sumram[94][133]+sumram[94][134]+sumram[94][135]+sumram[94][136];
    assign sumcache[95]=sumram[95][0]+sumram[95][1]+sumram[95][2]+sumram[95][3]+sumram[95][4]+sumram[95][5]+sumram[95][6]+sumram[95][7]+sumram[95][8]+sumram[95][9]+sumram[95][10]+sumram[95][11]+sumram[95][12]+sumram[95][13]+sumram[95][14]+sumram[95][15]+sumram[95][16]+sumram[95][17]+sumram[95][18]+sumram[95][19]+sumram[95][20]+sumram[95][21]+sumram[95][22]+sumram[95][23]+sumram[95][24]+sumram[95][25]+sumram[95][26]+sumram[95][27]+sumram[95][28]+sumram[95][29]+sumram[95][30]+sumram[95][31]+sumram[95][32]+sumram[95][33]+sumram[95][34]+sumram[95][35]+sumram[95][36]+sumram[95][37]+sumram[95][38]+sumram[95][39]+sumram[95][40]+sumram[95][41]+sumram[95][42]+sumram[95][43]+sumram[95][44]+sumram[95][45]+sumram[95][46]+sumram[95][47]+sumram[95][48]+sumram[95][49]+sumram[95][50]+sumram[95][51]+sumram[95][52]+sumram[95][53]+sumram[95][54]+sumram[95][55]+sumram[95][56]+sumram[95][57]+sumram[95][58]+sumram[95][59]+sumram[95][60]+sumram[95][61]+sumram[95][62]+sumram[95][63]+sumram[95][64]+sumram[95][65]+sumram[95][66]+sumram[95][67]+sumram[95][68]+sumram[95][69]+sumram[95][70]+sumram[95][71]+sumram[95][72]+sumram[95][73]+sumram[95][74]+sumram[95][75]+sumram[95][76]+sumram[95][77]+sumram[95][78]+sumram[95][79]+sumram[95][80]+sumram[95][81]+sumram[95][82]+sumram[95][83]+sumram[95][84]+sumram[95][85]+sumram[95][86]+sumram[95][87]+sumram[95][88]+sumram[95][89]+sumram[95][90]+sumram[95][91]+sumram[95][92]+sumram[95][93]+sumram[95][94]+sumram[95][95]+sumram[95][96]+sumram[95][97]+sumram[95][98]+sumram[95][99]+sumram[95][100]+sumram[95][101]+sumram[95][102]+sumram[95][103]+sumram[95][104]+sumram[95][105]+sumram[95][106]+sumram[95][107]+sumram[95][108]+sumram[95][109]+sumram[95][110]+sumram[95][111]+sumram[95][112]+sumram[95][113]+sumram[95][114]+sumram[95][115]+sumram[95][116]+sumram[95][117]+sumram[95][118]+sumram[95][119]+sumram[95][120]+sumram[95][121]+sumram[95][122]+sumram[95][123]+sumram[95][124]+sumram[95][125]+sumram[95][126]+sumram[95][127]+sumram[95][128]+sumram[95][129]+sumram[95][130]+sumram[95][131]+sumram[95][132]+sumram[95][133]+sumram[95][134]+sumram[95][135]+sumram[95][136];
    assign sumcache[96]=sumram[96][0]+sumram[96][1]+sumram[96][2]+sumram[96][3]+sumram[96][4]+sumram[96][5]+sumram[96][6]+sumram[96][7]+sumram[96][8]+sumram[96][9]+sumram[96][10]+sumram[96][11]+sumram[96][12]+sumram[96][13]+sumram[96][14]+sumram[96][15]+sumram[96][16]+sumram[96][17]+sumram[96][18]+sumram[96][19]+sumram[96][20]+sumram[96][21]+sumram[96][22]+sumram[96][23]+sumram[96][24]+sumram[96][25]+sumram[96][26]+sumram[96][27]+sumram[96][28]+sumram[96][29]+sumram[96][30]+sumram[96][31]+sumram[96][32]+sumram[96][33]+sumram[96][34]+sumram[96][35]+sumram[96][36]+sumram[96][37]+sumram[96][38]+sumram[96][39]+sumram[96][40]+sumram[96][41]+sumram[96][42]+sumram[96][43]+sumram[96][44]+sumram[96][45]+sumram[96][46]+sumram[96][47]+sumram[96][48]+sumram[96][49]+sumram[96][50]+sumram[96][51]+sumram[96][52]+sumram[96][53]+sumram[96][54]+sumram[96][55]+sumram[96][56]+sumram[96][57]+sumram[96][58]+sumram[96][59]+sumram[96][60]+sumram[96][61]+sumram[96][62]+sumram[96][63]+sumram[96][64]+sumram[96][65]+sumram[96][66]+sumram[96][67]+sumram[96][68]+sumram[96][69]+sumram[96][70]+sumram[96][71]+sumram[96][72]+sumram[96][73]+sumram[96][74]+sumram[96][75]+sumram[96][76]+sumram[96][77]+sumram[96][78]+sumram[96][79]+sumram[96][80]+sumram[96][81]+sumram[96][82]+sumram[96][83]+sumram[96][84]+sumram[96][85]+sumram[96][86]+sumram[96][87]+sumram[96][88]+sumram[96][89]+sumram[96][90]+sumram[96][91]+sumram[96][92]+sumram[96][93]+sumram[96][94]+sumram[96][95]+sumram[96][96]+sumram[96][97]+sumram[96][98]+sumram[96][99]+sumram[96][100]+sumram[96][101]+sumram[96][102]+sumram[96][103]+sumram[96][104]+sumram[96][105]+sumram[96][106]+sumram[96][107]+sumram[96][108]+sumram[96][109]+sumram[96][110]+sumram[96][111]+sumram[96][112]+sumram[96][113]+sumram[96][114]+sumram[96][115]+sumram[96][116]+sumram[96][117]+sumram[96][118]+sumram[96][119]+sumram[96][120]+sumram[96][121]+sumram[96][122]+sumram[96][123]+sumram[96][124]+sumram[96][125]+sumram[96][126]+sumram[96][127]+sumram[96][128]+sumram[96][129]+sumram[96][130]+sumram[96][131]+sumram[96][132]+sumram[96][133]+sumram[96][134]+sumram[96][135]+sumram[96][136];
    assign sumcache[97]=sumram[97][0]+sumram[97][1]+sumram[97][2]+sumram[97][3]+sumram[97][4]+sumram[97][5]+sumram[97][6]+sumram[97][7]+sumram[97][8]+sumram[97][9]+sumram[97][10]+sumram[97][11]+sumram[97][12]+sumram[97][13]+sumram[97][14]+sumram[97][15]+sumram[97][16]+sumram[97][17]+sumram[97][18]+sumram[97][19]+sumram[97][20]+sumram[97][21]+sumram[97][22]+sumram[97][23]+sumram[97][24]+sumram[97][25]+sumram[97][26]+sumram[97][27]+sumram[97][28]+sumram[97][29]+sumram[97][30]+sumram[97][31]+sumram[97][32]+sumram[97][33]+sumram[97][34]+sumram[97][35]+sumram[97][36]+sumram[97][37]+sumram[97][38]+sumram[97][39]+sumram[97][40]+sumram[97][41]+sumram[97][42]+sumram[97][43]+sumram[97][44]+sumram[97][45]+sumram[97][46]+sumram[97][47]+sumram[97][48]+sumram[97][49]+sumram[97][50]+sumram[97][51]+sumram[97][52]+sumram[97][53]+sumram[97][54]+sumram[97][55]+sumram[97][56]+sumram[97][57]+sumram[97][58]+sumram[97][59]+sumram[97][60]+sumram[97][61]+sumram[97][62]+sumram[97][63]+sumram[97][64]+sumram[97][65]+sumram[97][66]+sumram[97][67]+sumram[97][68]+sumram[97][69]+sumram[97][70]+sumram[97][71]+sumram[97][72]+sumram[97][73]+sumram[97][74]+sumram[97][75]+sumram[97][76]+sumram[97][77]+sumram[97][78]+sumram[97][79]+sumram[97][80]+sumram[97][81]+sumram[97][82]+sumram[97][83]+sumram[97][84]+sumram[97][85]+sumram[97][86]+sumram[97][87]+sumram[97][88]+sumram[97][89]+sumram[97][90]+sumram[97][91]+sumram[97][92]+sumram[97][93]+sumram[97][94]+sumram[97][95]+sumram[97][96]+sumram[97][97]+sumram[97][98]+sumram[97][99]+sumram[97][100]+sumram[97][101]+sumram[97][102]+sumram[97][103]+sumram[97][104]+sumram[97][105]+sumram[97][106]+sumram[97][107]+sumram[97][108]+sumram[97][109]+sumram[97][110]+sumram[97][111]+sumram[97][112]+sumram[97][113]+sumram[97][114]+sumram[97][115]+sumram[97][116]+sumram[97][117]+sumram[97][118]+sumram[97][119]+sumram[97][120]+sumram[97][121]+sumram[97][122]+sumram[97][123]+sumram[97][124]+sumram[97][125]+sumram[97][126]+sumram[97][127]+sumram[97][128]+sumram[97][129]+sumram[97][130]+sumram[97][131]+sumram[97][132]+sumram[97][133]+sumram[97][134]+sumram[97][135]+sumram[97][136];
    assign sumcache[98]=sumram[98][0]+sumram[98][1]+sumram[98][2]+sumram[98][3]+sumram[98][4]+sumram[98][5]+sumram[98][6]+sumram[98][7]+sumram[98][8]+sumram[98][9]+sumram[98][10]+sumram[98][11]+sumram[98][12]+sumram[98][13]+sumram[98][14]+sumram[98][15]+sumram[98][16]+sumram[98][17]+sumram[98][18]+sumram[98][19]+sumram[98][20]+sumram[98][21]+sumram[98][22]+sumram[98][23]+sumram[98][24]+sumram[98][25]+sumram[98][26]+sumram[98][27]+sumram[98][28]+sumram[98][29]+sumram[98][30]+sumram[98][31]+sumram[98][32]+sumram[98][33]+sumram[98][34]+sumram[98][35]+sumram[98][36]+sumram[98][37]+sumram[98][38]+sumram[98][39]+sumram[98][40]+sumram[98][41]+sumram[98][42]+sumram[98][43]+sumram[98][44]+sumram[98][45]+sumram[98][46]+sumram[98][47]+sumram[98][48]+sumram[98][49]+sumram[98][50]+sumram[98][51]+sumram[98][52]+sumram[98][53]+sumram[98][54]+sumram[98][55]+sumram[98][56]+sumram[98][57]+sumram[98][58]+sumram[98][59]+sumram[98][60]+sumram[98][61]+sumram[98][62]+sumram[98][63]+sumram[98][64]+sumram[98][65]+sumram[98][66]+sumram[98][67]+sumram[98][68]+sumram[98][69]+sumram[98][70]+sumram[98][71]+sumram[98][72]+sumram[98][73]+sumram[98][74]+sumram[98][75]+sumram[98][76]+sumram[98][77]+sumram[98][78]+sumram[98][79]+sumram[98][80]+sumram[98][81]+sumram[98][82]+sumram[98][83]+sumram[98][84]+sumram[98][85]+sumram[98][86]+sumram[98][87]+sumram[98][88]+sumram[98][89]+sumram[98][90]+sumram[98][91]+sumram[98][92]+sumram[98][93]+sumram[98][94]+sumram[98][95]+sumram[98][96]+sumram[98][97]+sumram[98][98]+sumram[98][99]+sumram[98][100]+sumram[98][101]+sumram[98][102]+sumram[98][103]+sumram[98][104]+sumram[98][105]+sumram[98][106]+sumram[98][107]+sumram[98][108]+sumram[98][109]+sumram[98][110]+sumram[98][111]+sumram[98][112]+sumram[98][113]+sumram[98][114]+sumram[98][115]+sumram[98][116]+sumram[98][117]+sumram[98][118]+sumram[98][119]+sumram[98][120]+sumram[98][121]+sumram[98][122]+sumram[98][123]+sumram[98][124]+sumram[98][125]+sumram[98][126]+sumram[98][127]+sumram[98][128]+sumram[98][129]+sumram[98][130]+sumram[98][131]+sumram[98][132]+sumram[98][133]+sumram[98][134]+sumram[98][135]+sumram[98][136];
    assign sumcache[99]=sumram[99][0]+sumram[99][1]+sumram[99][2]+sumram[99][3]+sumram[99][4]+sumram[99][5]+sumram[99][6]+sumram[99][7]+sumram[99][8]+sumram[99][9]+sumram[99][10]+sumram[99][11]+sumram[99][12]+sumram[99][13]+sumram[99][14]+sumram[99][15]+sumram[99][16]+sumram[99][17]+sumram[99][18]+sumram[99][19]+sumram[99][20]+sumram[99][21]+sumram[99][22]+sumram[99][23]+sumram[99][24]+sumram[99][25]+sumram[99][26]+sumram[99][27]+sumram[99][28]+sumram[99][29]+sumram[99][30]+sumram[99][31]+sumram[99][32]+sumram[99][33]+sumram[99][34]+sumram[99][35]+sumram[99][36]+sumram[99][37]+sumram[99][38]+sumram[99][39]+sumram[99][40]+sumram[99][41]+sumram[99][42]+sumram[99][43]+sumram[99][44]+sumram[99][45]+sumram[99][46]+sumram[99][47]+sumram[99][48]+sumram[99][49]+sumram[99][50]+sumram[99][51]+sumram[99][52]+sumram[99][53]+sumram[99][54]+sumram[99][55]+sumram[99][56]+sumram[99][57]+sumram[99][58]+sumram[99][59]+sumram[99][60]+sumram[99][61]+sumram[99][62]+sumram[99][63]+sumram[99][64]+sumram[99][65]+sumram[99][66]+sumram[99][67]+sumram[99][68]+sumram[99][69]+sumram[99][70]+sumram[99][71]+sumram[99][72]+sumram[99][73]+sumram[99][74]+sumram[99][75]+sumram[99][76]+sumram[99][77]+sumram[99][78]+sumram[99][79]+sumram[99][80]+sumram[99][81]+sumram[99][82]+sumram[99][83]+sumram[99][84]+sumram[99][85]+sumram[99][86]+sumram[99][87]+sumram[99][88]+sumram[99][89]+sumram[99][90]+sumram[99][91]+sumram[99][92]+sumram[99][93]+sumram[99][94]+sumram[99][95]+sumram[99][96]+sumram[99][97]+sumram[99][98]+sumram[99][99]+sumram[99][100]+sumram[99][101]+sumram[99][102]+sumram[99][103]+sumram[99][104]+sumram[99][105]+sumram[99][106]+sumram[99][107]+sumram[99][108]+sumram[99][109]+sumram[99][110]+sumram[99][111]+sumram[99][112]+sumram[99][113]+sumram[99][114]+sumram[99][115]+sumram[99][116]+sumram[99][117]+sumram[99][118]+sumram[99][119]+sumram[99][120]+sumram[99][121]+sumram[99][122]+sumram[99][123]+sumram[99][124]+sumram[99][125]+sumram[99][126]+sumram[99][127]+sumram[99][128]+sumram[99][129]+sumram[99][130]+sumram[99][131]+sumram[99][132]+sumram[99][133]+sumram[99][134]+sumram[99][135]+sumram[99][136];
    assign sumcache[100]=sumram[100][0]+sumram[100][1]+sumram[100][2]+sumram[100][3]+sumram[100][4]+sumram[100][5]+sumram[100][6]+sumram[100][7]+sumram[100][8]+sumram[100][9]+sumram[100][10]+sumram[100][11]+sumram[100][12]+sumram[100][13]+sumram[100][14]+sumram[100][15]+sumram[100][16]+sumram[100][17]+sumram[100][18]+sumram[100][19]+sumram[100][20]+sumram[100][21]+sumram[100][22]+sumram[100][23]+sumram[100][24]+sumram[100][25]+sumram[100][26]+sumram[100][27]+sumram[100][28]+sumram[100][29]+sumram[100][30]+sumram[100][31]+sumram[100][32]+sumram[100][33]+sumram[100][34]+sumram[100][35]+sumram[100][36]+sumram[100][37]+sumram[100][38]+sumram[100][39]+sumram[100][40]+sumram[100][41]+sumram[100][42]+sumram[100][43]+sumram[100][44]+sumram[100][45]+sumram[100][46]+sumram[100][47]+sumram[100][48]+sumram[100][49]+sumram[100][50]+sumram[100][51]+sumram[100][52]+sumram[100][53]+sumram[100][54]+sumram[100][55]+sumram[100][56]+sumram[100][57]+sumram[100][58]+sumram[100][59]+sumram[100][60]+sumram[100][61]+sumram[100][62]+sumram[100][63]+sumram[100][64]+sumram[100][65]+sumram[100][66]+sumram[100][67]+sumram[100][68]+sumram[100][69]+sumram[100][70]+sumram[100][71]+sumram[100][72]+sumram[100][73]+sumram[100][74]+sumram[100][75]+sumram[100][76]+sumram[100][77]+sumram[100][78]+sumram[100][79]+sumram[100][80]+sumram[100][81]+sumram[100][82]+sumram[100][83]+sumram[100][84]+sumram[100][85]+sumram[100][86]+sumram[100][87]+sumram[100][88]+sumram[100][89]+sumram[100][90]+sumram[100][91]+sumram[100][92]+sumram[100][93]+sumram[100][94]+sumram[100][95]+sumram[100][96]+sumram[100][97]+sumram[100][98]+sumram[100][99]+sumram[100][100]+sumram[100][101]+sumram[100][102]+sumram[100][103]+sumram[100][104]+sumram[100][105]+sumram[100][106]+sumram[100][107]+sumram[100][108]+sumram[100][109]+sumram[100][110]+sumram[100][111]+sumram[100][112]+sumram[100][113]+sumram[100][114]+sumram[100][115]+sumram[100][116]+sumram[100][117]+sumram[100][118]+sumram[100][119]+sumram[100][120]+sumram[100][121]+sumram[100][122]+sumram[100][123]+sumram[100][124]+sumram[100][125]+sumram[100][126]+sumram[100][127]+sumram[100][128]+sumram[100][129]+sumram[100][130]+sumram[100][131]+sumram[100][132]+sumram[100][133]+sumram[100][134]+sumram[100][135]+sumram[100][136];
    assign sumcache[101]=sumram[101][0]+sumram[101][1]+sumram[101][2]+sumram[101][3]+sumram[101][4]+sumram[101][5]+sumram[101][6]+sumram[101][7]+sumram[101][8]+sumram[101][9]+sumram[101][10]+sumram[101][11]+sumram[101][12]+sumram[101][13]+sumram[101][14]+sumram[101][15]+sumram[101][16]+sumram[101][17]+sumram[101][18]+sumram[101][19]+sumram[101][20]+sumram[101][21]+sumram[101][22]+sumram[101][23]+sumram[101][24]+sumram[101][25]+sumram[101][26]+sumram[101][27]+sumram[101][28]+sumram[101][29]+sumram[101][30]+sumram[101][31]+sumram[101][32]+sumram[101][33]+sumram[101][34]+sumram[101][35]+sumram[101][36]+sumram[101][37]+sumram[101][38]+sumram[101][39]+sumram[101][40]+sumram[101][41]+sumram[101][42]+sumram[101][43]+sumram[101][44]+sumram[101][45]+sumram[101][46]+sumram[101][47]+sumram[101][48]+sumram[101][49]+sumram[101][50]+sumram[101][51]+sumram[101][52]+sumram[101][53]+sumram[101][54]+sumram[101][55]+sumram[101][56]+sumram[101][57]+sumram[101][58]+sumram[101][59]+sumram[101][60]+sumram[101][61]+sumram[101][62]+sumram[101][63]+sumram[101][64]+sumram[101][65]+sumram[101][66]+sumram[101][67]+sumram[101][68]+sumram[101][69]+sumram[101][70]+sumram[101][71]+sumram[101][72]+sumram[101][73]+sumram[101][74]+sumram[101][75]+sumram[101][76]+sumram[101][77]+sumram[101][78]+sumram[101][79]+sumram[101][80]+sumram[101][81]+sumram[101][82]+sumram[101][83]+sumram[101][84]+sumram[101][85]+sumram[101][86]+sumram[101][87]+sumram[101][88]+sumram[101][89]+sumram[101][90]+sumram[101][91]+sumram[101][92]+sumram[101][93]+sumram[101][94]+sumram[101][95]+sumram[101][96]+sumram[101][97]+sumram[101][98]+sumram[101][99]+sumram[101][100]+sumram[101][101]+sumram[101][102]+sumram[101][103]+sumram[101][104]+sumram[101][105]+sumram[101][106]+sumram[101][107]+sumram[101][108]+sumram[101][109]+sumram[101][110]+sumram[101][111]+sumram[101][112]+sumram[101][113]+sumram[101][114]+sumram[101][115]+sumram[101][116]+sumram[101][117]+sumram[101][118]+sumram[101][119]+sumram[101][120]+sumram[101][121]+sumram[101][122]+sumram[101][123]+sumram[101][124]+sumram[101][125]+sumram[101][126]+sumram[101][127]+sumram[101][128]+sumram[101][129]+sumram[101][130]+sumram[101][131]+sumram[101][132]+sumram[101][133]+sumram[101][134]+sumram[101][135]+sumram[101][136];
    assign sumcache[102]=sumram[102][0]+sumram[102][1]+sumram[102][2]+sumram[102][3]+sumram[102][4]+sumram[102][5]+sumram[102][6]+sumram[102][7]+sumram[102][8]+sumram[102][9]+sumram[102][10]+sumram[102][11]+sumram[102][12]+sumram[102][13]+sumram[102][14]+sumram[102][15]+sumram[102][16]+sumram[102][17]+sumram[102][18]+sumram[102][19]+sumram[102][20]+sumram[102][21]+sumram[102][22]+sumram[102][23]+sumram[102][24]+sumram[102][25]+sumram[102][26]+sumram[102][27]+sumram[102][28]+sumram[102][29]+sumram[102][30]+sumram[102][31]+sumram[102][32]+sumram[102][33]+sumram[102][34]+sumram[102][35]+sumram[102][36]+sumram[102][37]+sumram[102][38]+sumram[102][39]+sumram[102][40]+sumram[102][41]+sumram[102][42]+sumram[102][43]+sumram[102][44]+sumram[102][45]+sumram[102][46]+sumram[102][47]+sumram[102][48]+sumram[102][49]+sumram[102][50]+sumram[102][51]+sumram[102][52]+sumram[102][53]+sumram[102][54]+sumram[102][55]+sumram[102][56]+sumram[102][57]+sumram[102][58]+sumram[102][59]+sumram[102][60]+sumram[102][61]+sumram[102][62]+sumram[102][63]+sumram[102][64]+sumram[102][65]+sumram[102][66]+sumram[102][67]+sumram[102][68]+sumram[102][69]+sumram[102][70]+sumram[102][71]+sumram[102][72]+sumram[102][73]+sumram[102][74]+sumram[102][75]+sumram[102][76]+sumram[102][77]+sumram[102][78]+sumram[102][79]+sumram[102][80]+sumram[102][81]+sumram[102][82]+sumram[102][83]+sumram[102][84]+sumram[102][85]+sumram[102][86]+sumram[102][87]+sumram[102][88]+sumram[102][89]+sumram[102][90]+sumram[102][91]+sumram[102][92]+sumram[102][93]+sumram[102][94]+sumram[102][95]+sumram[102][96]+sumram[102][97]+sumram[102][98]+sumram[102][99]+sumram[102][100]+sumram[102][101]+sumram[102][102]+sumram[102][103]+sumram[102][104]+sumram[102][105]+sumram[102][106]+sumram[102][107]+sumram[102][108]+sumram[102][109]+sumram[102][110]+sumram[102][111]+sumram[102][112]+sumram[102][113]+sumram[102][114]+sumram[102][115]+sumram[102][116]+sumram[102][117]+sumram[102][118]+sumram[102][119]+sumram[102][120]+sumram[102][121]+sumram[102][122]+sumram[102][123]+sumram[102][124]+sumram[102][125]+sumram[102][126]+sumram[102][127]+sumram[102][128]+sumram[102][129]+sumram[102][130]+sumram[102][131]+sumram[102][132]+sumram[102][133]+sumram[102][134]+sumram[102][135]+sumram[102][136];
    assign sumcache[103]=sumram[103][0]+sumram[103][1]+sumram[103][2]+sumram[103][3]+sumram[103][4]+sumram[103][5]+sumram[103][6]+sumram[103][7]+sumram[103][8]+sumram[103][9]+sumram[103][10]+sumram[103][11]+sumram[103][12]+sumram[103][13]+sumram[103][14]+sumram[103][15]+sumram[103][16]+sumram[103][17]+sumram[103][18]+sumram[103][19]+sumram[103][20]+sumram[103][21]+sumram[103][22]+sumram[103][23]+sumram[103][24]+sumram[103][25]+sumram[103][26]+sumram[103][27]+sumram[103][28]+sumram[103][29]+sumram[103][30]+sumram[103][31]+sumram[103][32]+sumram[103][33]+sumram[103][34]+sumram[103][35]+sumram[103][36]+sumram[103][37]+sumram[103][38]+sumram[103][39]+sumram[103][40]+sumram[103][41]+sumram[103][42]+sumram[103][43]+sumram[103][44]+sumram[103][45]+sumram[103][46]+sumram[103][47]+sumram[103][48]+sumram[103][49]+sumram[103][50]+sumram[103][51]+sumram[103][52]+sumram[103][53]+sumram[103][54]+sumram[103][55]+sumram[103][56]+sumram[103][57]+sumram[103][58]+sumram[103][59]+sumram[103][60]+sumram[103][61]+sumram[103][62]+sumram[103][63]+sumram[103][64]+sumram[103][65]+sumram[103][66]+sumram[103][67]+sumram[103][68]+sumram[103][69]+sumram[103][70]+sumram[103][71]+sumram[103][72]+sumram[103][73]+sumram[103][74]+sumram[103][75]+sumram[103][76]+sumram[103][77]+sumram[103][78]+sumram[103][79]+sumram[103][80]+sumram[103][81]+sumram[103][82]+sumram[103][83]+sumram[103][84]+sumram[103][85]+sumram[103][86]+sumram[103][87]+sumram[103][88]+sumram[103][89]+sumram[103][90]+sumram[103][91]+sumram[103][92]+sumram[103][93]+sumram[103][94]+sumram[103][95]+sumram[103][96]+sumram[103][97]+sumram[103][98]+sumram[103][99]+sumram[103][100]+sumram[103][101]+sumram[103][102]+sumram[103][103]+sumram[103][104]+sumram[103][105]+sumram[103][106]+sumram[103][107]+sumram[103][108]+sumram[103][109]+sumram[103][110]+sumram[103][111]+sumram[103][112]+sumram[103][113]+sumram[103][114]+sumram[103][115]+sumram[103][116]+sumram[103][117]+sumram[103][118]+sumram[103][119]+sumram[103][120]+sumram[103][121]+sumram[103][122]+sumram[103][123]+sumram[103][124]+sumram[103][125]+sumram[103][126]+sumram[103][127]+sumram[103][128]+sumram[103][129]+sumram[103][130]+sumram[103][131]+sumram[103][132]+sumram[103][133]+sumram[103][134]+sumram[103][135]+sumram[103][136];
    assign sumcache[104]=sumram[104][0]+sumram[104][1]+sumram[104][2]+sumram[104][3]+sumram[104][4]+sumram[104][5]+sumram[104][6]+sumram[104][7]+sumram[104][8]+sumram[104][9]+sumram[104][10]+sumram[104][11]+sumram[104][12]+sumram[104][13]+sumram[104][14]+sumram[104][15]+sumram[104][16]+sumram[104][17]+sumram[104][18]+sumram[104][19]+sumram[104][20]+sumram[104][21]+sumram[104][22]+sumram[104][23]+sumram[104][24]+sumram[104][25]+sumram[104][26]+sumram[104][27]+sumram[104][28]+sumram[104][29]+sumram[104][30]+sumram[104][31]+sumram[104][32]+sumram[104][33]+sumram[104][34]+sumram[104][35]+sumram[104][36]+sumram[104][37]+sumram[104][38]+sumram[104][39]+sumram[104][40]+sumram[104][41]+sumram[104][42]+sumram[104][43]+sumram[104][44]+sumram[104][45]+sumram[104][46]+sumram[104][47]+sumram[104][48]+sumram[104][49]+sumram[104][50]+sumram[104][51]+sumram[104][52]+sumram[104][53]+sumram[104][54]+sumram[104][55]+sumram[104][56]+sumram[104][57]+sumram[104][58]+sumram[104][59]+sumram[104][60]+sumram[104][61]+sumram[104][62]+sumram[104][63]+sumram[104][64]+sumram[104][65]+sumram[104][66]+sumram[104][67]+sumram[104][68]+sumram[104][69]+sumram[104][70]+sumram[104][71]+sumram[104][72]+sumram[104][73]+sumram[104][74]+sumram[104][75]+sumram[104][76]+sumram[104][77]+sumram[104][78]+sumram[104][79]+sumram[104][80]+sumram[104][81]+sumram[104][82]+sumram[104][83]+sumram[104][84]+sumram[104][85]+sumram[104][86]+sumram[104][87]+sumram[104][88]+sumram[104][89]+sumram[104][90]+sumram[104][91]+sumram[104][92]+sumram[104][93]+sumram[104][94]+sumram[104][95]+sumram[104][96]+sumram[104][97]+sumram[104][98]+sumram[104][99]+sumram[104][100]+sumram[104][101]+sumram[104][102]+sumram[104][103]+sumram[104][104]+sumram[104][105]+sumram[104][106]+sumram[104][107]+sumram[104][108]+sumram[104][109]+sumram[104][110]+sumram[104][111]+sumram[104][112]+sumram[104][113]+sumram[104][114]+sumram[104][115]+sumram[104][116]+sumram[104][117]+sumram[104][118]+sumram[104][119]+sumram[104][120]+sumram[104][121]+sumram[104][122]+sumram[104][123]+sumram[104][124]+sumram[104][125]+sumram[104][126]+sumram[104][127]+sumram[104][128]+sumram[104][129]+sumram[104][130]+sumram[104][131]+sumram[104][132]+sumram[104][133]+sumram[104][134]+sumram[104][135]+sumram[104][136];
    assign sumcache[105]=sumram[105][0]+sumram[105][1]+sumram[105][2]+sumram[105][3]+sumram[105][4]+sumram[105][5]+sumram[105][6]+sumram[105][7]+sumram[105][8]+sumram[105][9]+sumram[105][10]+sumram[105][11]+sumram[105][12]+sumram[105][13]+sumram[105][14]+sumram[105][15]+sumram[105][16]+sumram[105][17]+sumram[105][18]+sumram[105][19]+sumram[105][20]+sumram[105][21]+sumram[105][22]+sumram[105][23]+sumram[105][24]+sumram[105][25]+sumram[105][26]+sumram[105][27]+sumram[105][28]+sumram[105][29]+sumram[105][30]+sumram[105][31]+sumram[105][32]+sumram[105][33]+sumram[105][34]+sumram[105][35]+sumram[105][36]+sumram[105][37]+sumram[105][38]+sumram[105][39]+sumram[105][40]+sumram[105][41]+sumram[105][42]+sumram[105][43]+sumram[105][44]+sumram[105][45]+sumram[105][46]+sumram[105][47]+sumram[105][48]+sumram[105][49]+sumram[105][50]+sumram[105][51]+sumram[105][52]+sumram[105][53]+sumram[105][54]+sumram[105][55]+sumram[105][56]+sumram[105][57]+sumram[105][58]+sumram[105][59]+sumram[105][60]+sumram[105][61]+sumram[105][62]+sumram[105][63]+sumram[105][64]+sumram[105][65]+sumram[105][66]+sumram[105][67]+sumram[105][68]+sumram[105][69]+sumram[105][70]+sumram[105][71]+sumram[105][72]+sumram[105][73]+sumram[105][74]+sumram[105][75]+sumram[105][76]+sumram[105][77]+sumram[105][78]+sumram[105][79]+sumram[105][80]+sumram[105][81]+sumram[105][82]+sumram[105][83]+sumram[105][84]+sumram[105][85]+sumram[105][86]+sumram[105][87]+sumram[105][88]+sumram[105][89]+sumram[105][90]+sumram[105][91]+sumram[105][92]+sumram[105][93]+sumram[105][94]+sumram[105][95]+sumram[105][96]+sumram[105][97]+sumram[105][98]+sumram[105][99]+sumram[105][100]+sumram[105][101]+sumram[105][102]+sumram[105][103]+sumram[105][104]+sumram[105][105]+sumram[105][106]+sumram[105][107]+sumram[105][108]+sumram[105][109]+sumram[105][110]+sumram[105][111]+sumram[105][112]+sumram[105][113]+sumram[105][114]+sumram[105][115]+sumram[105][116]+sumram[105][117]+sumram[105][118]+sumram[105][119]+sumram[105][120]+sumram[105][121]+sumram[105][122]+sumram[105][123]+sumram[105][124]+sumram[105][125]+sumram[105][126]+sumram[105][127]+sumram[105][128]+sumram[105][129]+sumram[105][130]+sumram[105][131]+sumram[105][132]+sumram[105][133]+sumram[105][134]+sumram[105][135]+sumram[105][136];
    assign sumcache[106]=sumram[106][0]+sumram[106][1]+sumram[106][2]+sumram[106][3]+sumram[106][4]+sumram[106][5]+sumram[106][6]+sumram[106][7]+sumram[106][8]+sumram[106][9]+sumram[106][10]+sumram[106][11]+sumram[106][12]+sumram[106][13]+sumram[106][14]+sumram[106][15]+sumram[106][16]+sumram[106][17]+sumram[106][18]+sumram[106][19]+sumram[106][20]+sumram[106][21]+sumram[106][22]+sumram[106][23]+sumram[106][24]+sumram[106][25]+sumram[106][26]+sumram[106][27]+sumram[106][28]+sumram[106][29]+sumram[106][30]+sumram[106][31]+sumram[106][32]+sumram[106][33]+sumram[106][34]+sumram[106][35]+sumram[106][36]+sumram[106][37]+sumram[106][38]+sumram[106][39]+sumram[106][40]+sumram[106][41]+sumram[106][42]+sumram[106][43]+sumram[106][44]+sumram[106][45]+sumram[106][46]+sumram[106][47]+sumram[106][48]+sumram[106][49]+sumram[106][50]+sumram[106][51]+sumram[106][52]+sumram[106][53]+sumram[106][54]+sumram[106][55]+sumram[106][56]+sumram[106][57]+sumram[106][58]+sumram[106][59]+sumram[106][60]+sumram[106][61]+sumram[106][62]+sumram[106][63]+sumram[106][64]+sumram[106][65]+sumram[106][66]+sumram[106][67]+sumram[106][68]+sumram[106][69]+sumram[106][70]+sumram[106][71]+sumram[106][72]+sumram[106][73]+sumram[106][74]+sumram[106][75]+sumram[106][76]+sumram[106][77]+sumram[106][78]+sumram[106][79]+sumram[106][80]+sumram[106][81]+sumram[106][82]+sumram[106][83]+sumram[106][84]+sumram[106][85]+sumram[106][86]+sumram[106][87]+sumram[106][88]+sumram[106][89]+sumram[106][90]+sumram[106][91]+sumram[106][92]+sumram[106][93]+sumram[106][94]+sumram[106][95]+sumram[106][96]+sumram[106][97]+sumram[106][98]+sumram[106][99]+sumram[106][100]+sumram[106][101]+sumram[106][102]+sumram[106][103]+sumram[106][104]+sumram[106][105]+sumram[106][106]+sumram[106][107]+sumram[106][108]+sumram[106][109]+sumram[106][110]+sumram[106][111]+sumram[106][112]+sumram[106][113]+sumram[106][114]+sumram[106][115]+sumram[106][116]+sumram[106][117]+sumram[106][118]+sumram[106][119]+sumram[106][120]+sumram[106][121]+sumram[106][122]+sumram[106][123]+sumram[106][124]+sumram[106][125]+sumram[106][126]+sumram[106][127]+sumram[106][128]+sumram[106][129]+sumram[106][130]+sumram[106][131]+sumram[106][132]+sumram[106][133]+sumram[106][134]+sumram[106][135]+sumram[106][136];
    assign sumcache[107]=sumram[107][0]+sumram[107][1]+sumram[107][2]+sumram[107][3]+sumram[107][4]+sumram[107][5]+sumram[107][6]+sumram[107][7]+sumram[107][8]+sumram[107][9]+sumram[107][10]+sumram[107][11]+sumram[107][12]+sumram[107][13]+sumram[107][14]+sumram[107][15]+sumram[107][16]+sumram[107][17]+sumram[107][18]+sumram[107][19]+sumram[107][20]+sumram[107][21]+sumram[107][22]+sumram[107][23]+sumram[107][24]+sumram[107][25]+sumram[107][26]+sumram[107][27]+sumram[107][28]+sumram[107][29]+sumram[107][30]+sumram[107][31]+sumram[107][32]+sumram[107][33]+sumram[107][34]+sumram[107][35]+sumram[107][36]+sumram[107][37]+sumram[107][38]+sumram[107][39]+sumram[107][40]+sumram[107][41]+sumram[107][42]+sumram[107][43]+sumram[107][44]+sumram[107][45]+sumram[107][46]+sumram[107][47]+sumram[107][48]+sumram[107][49]+sumram[107][50]+sumram[107][51]+sumram[107][52]+sumram[107][53]+sumram[107][54]+sumram[107][55]+sumram[107][56]+sumram[107][57]+sumram[107][58]+sumram[107][59]+sumram[107][60]+sumram[107][61]+sumram[107][62]+sumram[107][63]+sumram[107][64]+sumram[107][65]+sumram[107][66]+sumram[107][67]+sumram[107][68]+sumram[107][69]+sumram[107][70]+sumram[107][71]+sumram[107][72]+sumram[107][73]+sumram[107][74]+sumram[107][75]+sumram[107][76]+sumram[107][77]+sumram[107][78]+sumram[107][79]+sumram[107][80]+sumram[107][81]+sumram[107][82]+sumram[107][83]+sumram[107][84]+sumram[107][85]+sumram[107][86]+sumram[107][87]+sumram[107][88]+sumram[107][89]+sumram[107][90]+sumram[107][91]+sumram[107][92]+sumram[107][93]+sumram[107][94]+sumram[107][95]+sumram[107][96]+sumram[107][97]+sumram[107][98]+sumram[107][99]+sumram[107][100]+sumram[107][101]+sumram[107][102]+sumram[107][103]+sumram[107][104]+sumram[107][105]+sumram[107][106]+sumram[107][107]+sumram[107][108]+sumram[107][109]+sumram[107][110]+sumram[107][111]+sumram[107][112]+sumram[107][113]+sumram[107][114]+sumram[107][115]+sumram[107][116]+sumram[107][117]+sumram[107][118]+sumram[107][119]+sumram[107][120]+sumram[107][121]+sumram[107][122]+sumram[107][123]+sumram[107][124]+sumram[107][125]+sumram[107][126]+sumram[107][127]+sumram[107][128]+sumram[107][129]+sumram[107][130]+sumram[107][131]+sumram[107][132]+sumram[107][133]+sumram[107][134]+sumram[107][135]+sumram[107][136];
    assign sumcache[108]=sumram[108][0]+sumram[108][1]+sumram[108][2]+sumram[108][3]+sumram[108][4]+sumram[108][5]+sumram[108][6]+sumram[108][7]+sumram[108][8]+sumram[108][9]+sumram[108][10]+sumram[108][11]+sumram[108][12]+sumram[108][13]+sumram[108][14]+sumram[108][15]+sumram[108][16]+sumram[108][17]+sumram[108][18]+sumram[108][19]+sumram[108][20]+sumram[108][21]+sumram[108][22]+sumram[108][23]+sumram[108][24]+sumram[108][25]+sumram[108][26]+sumram[108][27]+sumram[108][28]+sumram[108][29]+sumram[108][30]+sumram[108][31]+sumram[108][32]+sumram[108][33]+sumram[108][34]+sumram[108][35]+sumram[108][36]+sumram[108][37]+sumram[108][38]+sumram[108][39]+sumram[108][40]+sumram[108][41]+sumram[108][42]+sumram[108][43]+sumram[108][44]+sumram[108][45]+sumram[108][46]+sumram[108][47]+sumram[108][48]+sumram[108][49]+sumram[108][50]+sumram[108][51]+sumram[108][52]+sumram[108][53]+sumram[108][54]+sumram[108][55]+sumram[108][56]+sumram[108][57]+sumram[108][58]+sumram[108][59]+sumram[108][60]+sumram[108][61]+sumram[108][62]+sumram[108][63]+sumram[108][64]+sumram[108][65]+sumram[108][66]+sumram[108][67]+sumram[108][68]+sumram[108][69]+sumram[108][70]+sumram[108][71]+sumram[108][72]+sumram[108][73]+sumram[108][74]+sumram[108][75]+sumram[108][76]+sumram[108][77]+sumram[108][78]+sumram[108][79]+sumram[108][80]+sumram[108][81]+sumram[108][82]+sumram[108][83]+sumram[108][84]+sumram[108][85]+sumram[108][86]+sumram[108][87]+sumram[108][88]+sumram[108][89]+sumram[108][90]+sumram[108][91]+sumram[108][92]+sumram[108][93]+sumram[108][94]+sumram[108][95]+sumram[108][96]+sumram[108][97]+sumram[108][98]+sumram[108][99]+sumram[108][100]+sumram[108][101]+sumram[108][102]+sumram[108][103]+sumram[108][104]+sumram[108][105]+sumram[108][106]+sumram[108][107]+sumram[108][108]+sumram[108][109]+sumram[108][110]+sumram[108][111]+sumram[108][112]+sumram[108][113]+sumram[108][114]+sumram[108][115]+sumram[108][116]+sumram[108][117]+sumram[108][118]+sumram[108][119]+sumram[108][120]+sumram[108][121]+sumram[108][122]+sumram[108][123]+sumram[108][124]+sumram[108][125]+sumram[108][126]+sumram[108][127]+sumram[108][128]+sumram[108][129]+sumram[108][130]+sumram[108][131]+sumram[108][132]+sumram[108][133]+sumram[108][134]+sumram[108][135]+sumram[108][136];
    assign sumcache[109]=sumram[109][0]+sumram[109][1]+sumram[109][2]+sumram[109][3]+sumram[109][4]+sumram[109][5]+sumram[109][6]+sumram[109][7]+sumram[109][8]+sumram[109][9]+sumram[109][10]+sumram[109][11]+sumram[109][12]+sumram[109][13]+sumram[109][14]+sumram[109][15]+sumram[109][16]+sumram[109][17]+sumram[109][18]+sumram[109][19]+sumram[109][20]+sumram[109][21]+sumram[109][22]+sumram[109][23]+sumram[109][24]+sumram[109][25]+sumram[109][26]+sumram[109][27]+sumram[109][28]+sumram[109][29]+sumram[109][30]+sumram[109][31]+sumram[109][32]+sumram[109][33]+sumram[109][34]+sumram[109][35]+sumram[109][36]+sumram[109][37]+sumram[109][38]+sumram[109][39]+sumram[109][40]+sumram[109][41]+sumram[109][42]+sumram[109][43]+sumram[109][44]+sumram[109][45]+sumram[109][46]+sumram[109][47]+sumram[109][48]+sumram[109][49]+sumram[109][50]+sumram[109][51]+sumram[109][52]+sumram[109][53]+sumram[109][54]+sumram[109][55]+sumram[109][56]+sumram[109][57]+sumram[109][58]+sumram[109][59]+sumram[109][60]+sumram[109][61]+sumram[109][62]+sumram[109][63]+sumram[109][64]+sumram[109][65]+sumram[109][66]+sumram[109][67]+sumram[109][68]+sumram[109][69]+sumram[109][70]+sumram[109][71]+sumram[109][72]+sumram[109][73]+sumram[109][74]+sumram[109][75]+sumram[109][76]+sumram[109][77]+sumram[109][78]+sumram[109][79]+sumram[109][80]+sumram[109][81]+sumram[109][82]+sumram[109][83]+sumram[109][84]+sumram[109][85]+sumram[109][86]+sumram[109][87]+sumram[109][88]+sumram[109][89]+sumram[109][90]+sumram[109][91]+sumram[109][92]+sumram[109][93]+sumram[109][94]+sumram[109][95]+sumram[109][96]+sumram[109][97]+sumram[109][98]+sumram[109][99]+sumram[109][100]+sumram[109][101]+sumram[109][102]+sumram[109][103]+sumram[109][104]+sumram[109][105]+sumram[109][106]+sumram[109][107]+sumram[109][108]+sumram[109][109]+sumram[109][110]+sumram[109][111]+sumram[109][112]+sumram[109][113]+sumram[109][114]+sumram[109][115]+sumram[109][116]+sumram[109][117]+sumram[109][118]+sumram[109][119]+sumram[109][120]+sumram[109][121]+sumram[109][122]+sumram[109][123]+sumram[109][124]+sumram[109][125]+sumram[109][126]+sumram[109][127]+sumram[109][128]+sumram[109][129]+sumram[109][130]+sumram[109][131]+sumram[109][132]+sumram[109][133]+sumram[109][134]+sumram[109][135]+sumram[109][136];
    assign sumcache[110]=sumram[110][0]+sumram[110][1]+sumram[110][2]+sumram[110][3]+sumram[110][4]+sumram[110][5]+sumram[110][6]+sumram[110][7]+sumram[110][8]+sumram[110][9]+sumram[110][10]+sumram[110][11]+sumram[110][12]+sumram[110][13]+sumram[110][14]+sumram[110][15]+sumram[110][16]+sumram[110][17]+sumram[110][18]+sumram[110][19]+sumram[110][20]+sumram[110][21]+sumram[110][22]+sumram[110][23]+sumram[110][24]+sumram[110][25]+sumram[110][26]+sumram[110][27]+sumram[110][28]+sumram[110][29]+sumram[110][30]+sumram[110][31]+sumram[110][32]+sumram[110][33]+sumram[110][34]+sumram[110][35]+sumram[110][36]+sumram[110][37]+sumram[110][38]+sumram[110][39]+sumram[110][40]+sumram[110][41]+sumram[110][42]+sumram[110][43]+sumram[110][44]+sumram[110][45]+sumram[110][46]+sumram[110][47]+sumram[110][48]+sumram[110][49]+sumram[110][50]+sumram[110][51]+sumram[110][52]+sumram[110][53]+sumram[110][54]+sumram[110][55]+sumram[110][56]+sumram[110][57]+sumram[110][58]+sumram[110][59]+sumram[110][60]+sumram[110][61]+sumram[110][62]+sumram[110][63]+sumram[110][64]+sumram[110][65]+sumram[110][66]+sumram[110][67]+sumram[110][68]+sumram[110][69]+sumram[110][70]+sumram[110][71]+sumram[110][72]+sumram[110][73]+sumram[110][74]+sumram[110][75]+sumram[110][76]+sumram[110][77]+sumram[110][78]+sumram[110][79]+sumram[110][80]+sumram[110][81]+sumram[110][82]+sumram[110][83]+sumram[110][84]+sumram[110][85]+sumram[110][86]+sumram[110][87]+sumram[110][88]+sumram[110][89]+sumram[110][90]+sumram[110][91]+sumram[110][92]+sumram[110][93]+sumram[110][94]+sumram[110][95]+sumram[110][96]+sumram[110][97]+sumram[110][98]+sumram[110][99]+sumram[110][100]+sumram[110][101]+sumram[110][102]+sumram[110][103]+sumram[110][104]+sumram[110][105]+sumram[110][106]+sumram[110][107]+sumram[110][108]+sumram[110][109]+sumram[110][110]+sumram[110][111]+sumram[110][112]+sumram[110][113]+sumram[110][114]+sumram[110][115]+sumram[110][116]+sumram[110][117]+sumram[110][118]+sumram[110][119]+sumram[110][120]+sumram[110][121]+sumram[110][122]+sumram[110][123]+sumram[110][124]+sumram[110][125]+sumram[110][126]+sumram[110][127]+sumram[110][128]+sumram[110][129]+sumram[110][130]+sumram[110][131]+sumram[110][132]+sumram[110][133]+sumram[110][134]+sumram[110][135]+sumram[110][136];
    assign sumcache[111]=sumram[111][0]+sumram[111][1]+sumram[111][2]+sumram[111][3]+sumram[111][4]+sumram[111][5]+sumram[111][6]+sumram[111][7]+sumram[111][8]+sumram[111][9]+sumram[111][10]+sumram[111][11]+sumram[111][12]+sumram[111][13]+sumram[111][14]+sumram[111][15]+sumram[111][16]+sumram[111][17]+sumram[111][18]+sumram[111][19]+sumram[111][20]+sumram[111][21]+sumram[111][22]+sumram[111][23]+sumram[111][24]+sumram[111][25]+sumram[111][26]+sumram[111][27]+sumram[111][28]+sumram[111][29]+sumram[111][30]+sumram[111][31]+sumram[111][32]+sumram[111][33]+sumram[111][34]+sumram[111][35]+sumram[111][36]+sumram[111][37]+sumram[111][38]+sumram[111][39]+sumram[111][40]+sumram[111][41]+sumram[111][42]+sumram[111][43]+sumram[111][44]+sumram[111][45]+sumram[111][46]+sumram[111][47]+sumram[111][48]+sumram[111][49]+sumram[111][50]+sumram[111][51]+sumram[111][52]+sumram[111][53]+sumram[111][54]+sumram[111][55]+sumram[111][56]+sumram[111][57]+sumram[111][58]+sumram[111][59]+sumram[111][60]+sumram[111][61]+sumram[111][62]+sumram[111][63]+sumram[111][64]+sumram[111][65]+sumram[111][66]+sumram[111][67]+sumram[111][68]+sumram[111][69]+sumram[111][70]+sumram[111][71]+sumram[111][72]+sumram[111][73]+sumram[111][74]+sumram[111][75]+sumram[111][76]+sumram[111][77]+sumram[111][78]+sumram[111][79]+sumram[111][80]+sumram[111][81]+sumram[111][82]+sumram[111][83]+sumram[111][84]+sumram[111][85]+sumram[111][86]+sumram[111][87]+sumram[111][88]+sumram[111][89]+sumram[111][90]+sumram[111][91]+sumram[111][92]+sumram[111][93]+sumram[111][94]+sumram[111][95]+sumram[111][96]+sumram[111][97]+sumram[111][98]+sumram[111][99]+sumram[111][100]+sumram[111][101]+sumram[111][102]+sumram[111][103]+sumram[111][104]+sumram[111][105]+sumram[111][106]+sumram[111][107]+sumram[111][108]+sumram[111][109]+sumram[111][110]+sumram[111][111]+sumram[111][112]+sumram[111][113]+sumram[111][114]+sumram[111][115]+sumram[111][116]+sumram[111][117]+sumram[111][118]+sumram[111][119]+sumram[111][120]+sumram[111][121]+sumram[111][122]+sumram[111][123]+sumram[111][124]+sumram[111][125]+sumram[111][126]+sumram[111][127]+sumram[111][128]+sumram[111][129]+sumram[111][130]+sumram[111][131]+sumram[111][132]+sumram[111][133]+sumram[111][134]+sumram[111][135]+sumram[111][136];
    assign sumcache[112]=sumram[112][0]+sumram[112][1]+sumram[112][2]+sumram[112][3]+sumram[112][4]+sumram[112][5]+sumram[112][6]+sumram[112][7]+sumram[112][8]+sumram[112][9]+sumram[112][10]+sumram[112][11]+sumram[112][12]+sumram[112][13]+sumram[112][14]+sumram[112][15]+sumram[112][16]+sumram[112][17]+sumram[112][18]+sumram[112][19]+sumram[112][20]+sumram[112][21]+sumram[112][22]+sumram[112][23]+sumram[112][24]+sumram[112][25]+sumram[112][26]+sumram[112][27]+sumram[112][28]+sumram[112][29]+sumram[112][30]+sumram[112][31]+sumram[112][32]+sumram[112][33]+sumram[112][34]+sumram[112][35]+sumram[112][36]+sumram[112][37]+sumram[112][38]+sumram[112][39]+sumram[112][40]+sumram[112][41]+sumram[112][42]+sumram[112][43]+sumram[112][44]+sumram[112][45]+sumram[112][46]+sumram[112][47]+sumram[112][48]+sumram[112][49]+sumram[112][50]+sumram[112][51]+sumram[112][52]+sumram[112][53]+sumram[112][54]+sumram[112][55]+sumram[112][56]+sumram[112][57]+sumram[112][58]+sumram[112][59]+sumram[112][60]+sumram[112][61]+sumram[112][62]+sumram[112][63]+sumram[112][64]+sumram[112][65]+sumram[112][66]+sumram[112][67]+sumram[112][68]+sumram[112][69]+sumram[112][70]+sumram[112][71]+sumram[112][72]+sumram[112][73]+sumram[112][74]+sumram[112][75]+sumram[112][76]+sumram[112][77]+sumram[112][78]+sumram[112][79]+sumram[112][80]+sumram[112][81]+sumram[112][82]+sumram[112][83]+sumram[112][84]+sumram[112][85]+sumram[112][86]+sumram[112][87]+sumram[112][88]+sumram[112][89]+sumram[112][90]+sumram[112][91]+sumram[112][92]+sumram[112][93]+sumram[112][94]+sumram[112][95]+sumram[112][96]+sumram[112][97]+sumram[112][98]+sumram[112][99]+sumram[112][100]+sumram[112][101]+sumram[112][102]+sumram[112][103]+sumram[112][104]+sumram[112][105]+sumram[112][106]+sumram[112][107]+sumram[112][108]+sumram[112][109]+sumram[112][110]+sumram[112][111]+sumram[112][112]+sumram[112][113]+sumram[112][114]+sumram[112][115]+sumram[112][116]+sumram[112][117]+sumram[112][118]+sumram[112][119]+sumram[112][120]+sumram[112][121]+sumram[112][122]+sumram[112][123]+sumram[112][124]+sumram[112][125]+sumram[112][126]+sumram[112][127]+sumram[112][128]+sumram[112][129]+sumram[112][130]+sumram[112][131]+sumram[112][132]+sumram[112][133]+sumram[112][134]+sumram[112][135]+sumram[112][136];
    assign sumcache[113]=sumram[113][0]+sumram[113][1]+sumram[113][2]+sumram[113][3]+sumram[113][4]+sumram[113][5]+sumram[113][6]+sumram[113][7]+sumram[113][8]+sumram[113][9]+sumram[113][10]+sumram[113][11]+sumram[113][12]+sumram[113][13]+sumram[113][14]+sumram[113][15]+sumram[113][16]+sumram[113][17]+sumram[113][18]+sumram[113][19]+sumram[113][20]+sumram[113][21]+sumram[113][22]+sumram[113][23]+sumram[113][24]+sumram[113][25]+sumram[113][26]+sumram[113][27]+sumram[113][28]+sumram[113][29]+sumram[113][30]+sumram[113][31]+sumram[113][32]+sumram[113][33]+sumram[113][34]+sumram[113][35]+sumram[113][36]+sumram[113][37]+sumram[113][38]+sumram[113][39]+sumram[113][40]+sumram[113][41]+sumram[113][42]+sumram[113][43]+sumram[113][44]+sumram[113][45]+sumram[113][46]+sumram[113][47]+sumram[113][48]+sumram[113][49]+sumram[113][50]+sumram[113][51]+sumram[113][52]+sumram[113][53]+sumram[113][54]+sumram[113][55]+sumram[113][56]+sumram[113][57]+sumram[113][58]+sumram[113][59]+sumram[113][60]+sumram[113][61]+sumram[113][62]+sumram[113][63]+sumram[113][64]+sumram[113][65]+sumram[113][66]+sumram[113][67]+sumram[113][68]+sumram[113][69]+sumram[113][70]+sumram[113][71]+sumram[113][72]+sumram[113][73]+sumram[113][74]+sumram[113][75]+sumram[113][76]+sumram[113][77]+sumram[113][78]+sumram[113][79]+sumram[113][80]+sumram[113][81]+sumram[113][82]+sumram[113][83]+sumram[113][84]+sumram[113][85]+sumram[113][86]+sumram[113][87]+sumram[113][88]+sumram[113][89]+sumram[113][90]+sumram[113][91]+sumram[113][92]+sumram[113][93]+sumram[113][94]+sumram[113][95]+sumram[113][96]+sumram[113][97]+sumram[113][98]+sumram[113][99]+sumram[113][100]+sumram[113][101]+sumram[113][102]+sumram[113][103]+sumram[113][104]+sumram[113][105]+sumram[113][106]+sumram[113][107]+sumram[113][108]+sumram[113][109]+sumram[113][110]+sumram[113][111]+sumram[113][112]+sumram[113][113]+sumram[113][114]+sumram[113][115]+sumram[113][116]+sumram[113][117]+sumram[113][118]+sumram[113][119]+sumram[113][120]+sumram[113][121]+sumram[113][122]+sumram[113][123]+sumram[113][124]+sumram[113][125]+sumram[113][126]+sumram[113][127]+sumram[113][128]+sumram[113][129]+sumram[113][130]+sumram[113][131]+sumram[113][132]+sumram[113][133]+sumram[113][134]+sumram[113][135]+sumram[113][136];
    assign sumcache[114]=sumram[114][0]+sumram[114][1]+sumram[114][2]+sumram[114][3]+sumram[114][4]+sumram[114][5]+sumram[114][6]+sumram[114][7]+sumram[114][8]+sumram[114][9]+sumram[114][10]+sumram[114][11]+sumram[114][12]+sumram[114][13]+sumram[114][14]+sumram[114][15]+sumram[114][16]+sumram[114][17]+sumram[114][18]+sumram[114][19]+sumram[114][20]+sumram[114][21]+sumram[114][22]+sumram[114][23]+sumram[114][24]+sumram[114][25]+sumram[114][26]+sumram[114][27]+sumram[114][28]+sumram[114][29]+sumram[114][30]+sumram[114][31]+sumram[114][32]+sumram[114][33]+sumram[114][34]+sumram[114][35]+sumram[114][36]+sumram[114][37]+sumram[114][38]+sumram[114][39]+sumram[114][40]+sumram[114][41]+sumram[114][42]+sumram[114][43]+sumram[114][44]+sumram[114][45]+sumram[114][46]+sumram[114][47]+sumram[114][48]+sumram[114][49]+sumram[114][50]+sumram[114][51]+sumram[114][52]+sumram[114][53]+sumram[114][54]+sumram[114][55]+sumram[114][56]+sumram[114][57]+sumram[114][58]+sumram[114][59]+sumram[114][60]+sumram[114][61]+sumram[114][62]+sumram[114][63]+sumram[114][64]+sumram[114][65]+sumram[114][66]+sumram[114][67]+sumram[114][68]+sumram[114][69]+sumram[114][70]+sumram[114][71]+sumram[114][72]+sumram[114][73]+sumram[114][74]+sumram[114][75]+sumram[114][76]+sumram[114][77]+sumram[114][78]+sumram[114][79]+sumram[114][80]+sumram[114][81]+sumram[114][82]+sumram[114][83]+sumram[114][84]+sumram[114][85]+sumram[114][86]+sumram[114][87]+sumram[114][88]+sumram[114][89]+sumram[114][90]+sumram[114][91]+sumram[114][92]+sumram[114][93]+sumram[114][94]+sumram[114][95]+sumram[114][96]+sumram[114][97]+sumram[114][98]+sumram[114][99]+sumram[114][100]+sumram[114][101]+sumram[114][102]+sumram[114][103]+sumram[114][104]+sumram[114][105]+sumram[114][106]+sumram[114][107]+sumram[114][108]+sumram[114][109]+sumram[114][110]+sumram[114][111]+sumram[114][112]+sumram[114][113]+sumram[114][114]+sumram[114][115]+sumram[114][116]+sumram[114][117]+sumram[114][118]+sumram[114][119]+sumram[114][120]+sumram[114][121]+sumram[114][122]+sumram[114][123]+sumram[114][124]+sumram[114][125]+sumram[114][126]+sumram[114][127]+sumram[114][128]+sumram[114][129]+sumram[114][130]+sumram[114][131]+sumram[114][132]+sumram[114][133]+sumram[114][134]+sumram[114][135]+sumram[114][136];
    assign sumcache[115]=sumram[115][0]+sumram[115][1]+sumram[115][2]+sumram[115][3]+sumram[115][4]+sumram[115][5]+sumram[115][6]+sumram[115][7]+sumram[115][8]+sumram[115][9]+sumram[115][10]+sumram[115][11]+sumram[115][12]+sumram[115][13]+sumram[115][14]+sumram[115][15]+sumram[115][16]+sumram[115][17]+sumram[115][18]+sumram[115][19]+sumram[115][20]+sumram[115][21]+sumram[115][22]+sumram[115][23]+sumram[115][24]+sumram[115][25]+sumram[115][26]+sumram[115][27]+sumram[115][28]+sumram[115][29]+sumram[115][30]+sumram[115][31]+sumram[115][32]+sumram[115][33]+sumram[115][34]+sumram[115][35]+sumram[115][36]+sumram[115][37]+sumram[115][38]+sumram[115][39]+sumram[115][40]+sumram[115][41]+sumram[115][42]+sumram[115][43]+sumram[115][44]+sumram[115][45]+sumram[115][46]+sumram[115][47]+sumram[115][48]+sumram[115][49]+sumram[115][50]+sumram[115][51]+sumram[115][52]+sumram[115][53]+sumram[115][54]+sumram[115][55]+sumram[115][56]+sumram[115][57]+sumram[115][58]+sumram[115][59]+sumram[115][60]+sumram[115][61]+sumram[115][62]+sumram[115][63]+sumram[115][64]+sumram[115][65]+sumram[115][66]+sumram[115][67]+sumram[115][68]+sumram[115][69]+sumram[115][70]+sumram[115][71]+sumram[115][72]+sumram[115][73]+sumram[115][74]+sumram[115][75]+sumram[115][76]+sumram[115][77]+sumram[115][78]+sumram[115][79]+sumram[115][80]+sumram[115][81]+sumram[115][82]+sumram[115][83]+sumram[115][84]+sumram[115][85]+sumram[115][86]+sumram[115][87]+sumram[115][88]+sumram[115][89]+sumram[115][90]+sumram[115][91]+sumram[115][92]+sumram[115][93]+sumram[115][94]+sumram[115][95]+sumram[115][96]+sumram[115][97]+sumram[115][98]+sumram[115][99]+sumram[115][100]+sumram[115][101]+sumram[115][102]+sumram[115][103]+sumram[115][104]+sumram[115][105]+sumram[115][106]+sumram[115][107]+sumram[115][108]+sumram[115][109]+sumram[115][110]+sumram[115][111]+sumram[115][112]+sumram[115][113]+sumram[115][114]+sumram[115][115]+sumram[115][116]+sumram[115][117]+sumram[115][118]+sumram[115][119]+sumram[115][120]+sumram[115][121]+sumram[115][122]+sumram[115][123]+sumram[115][124]+sumram[115][125]+sumram[115][126]+sumram[115][127]+sumram[115][128]+sumram[115][129]+sumram[115][130]+sumram[115][131]+sumram[115][132]+sumram[115][133]+sumram[115][134]+sumram[115][135]+sumram[115][136];
    assign sumcache[116]=sumram[116][0]+sumram[116][1]+sumram[116][2]+sumram[116][3]+sumram[116][4]+sumram[116][5]+sumram[116][6]+sumram[116][7]+sumram[116][8]+sumram[116][9]+sumram[116][10]+sumram[116][11]+sumram[116][12]+sumram[116][13]+sumram[116][14]+sumram[116][15]+sumram[116][16]+sumram[116][17]+sumram[116][18]+sumram[116][19]+sumram[116][20]+sumram[116][21]+sumram[116][22]+sumram[116][23]+sumram[116][24]+sumram[116][25]+sumram[116][26]+sumram[116][27]+sumram[116][28]+sumram[116][29]+sumram[116][30]+sumram[116][31]+sumram[116][32]+sumram[116][33]+sumram[116][34]+sumram[116][35]+sumram[116][36]+sumram[116][37]+sumram[116][38]+sumram[116][39]+sumram[116][40]+sumram[116][41]+sumram[116][42]+sumram[116][43]+sumram[116][44]+sumram[116][45]+sumram[116][46]+sumram[116][47]+sumram[116][48]+sumram[116][49]+sumram[116][50]+sumram[116][51]+sumram[116][52]+sumram[116][53]+sumram[116][54]+sumram[116][55]+sumram[116][56]+sumram[116][57]+sumram[116][58]+sumram[116][59]+sumram[116][60]+sumram[116][61]+sumram[116][62]+sumram[116][63]+sumram[116][64]+sumram[116][65]+sumram[116][66]+sumram[116][67]+sumram[116][68]+sumram[116][69]+sumram[116][70]+sumram[116][71]+sumram[116][72]+sumram[116][73]+sumram[116][74]+sumram[116][75]+sumram[116][76]+sumram[116][77]+sumram[116][78]+sumram[116][79]+sumram[116][80]+sumram[116][81]+sumram[116][82]+sumram[116][83]+sumram[116][84]+sumram[116][85]+sumram[116][86]+sumram[116][87]+sumram[116][88]+sumram[116][89]+sumram[116][90]+sumram[116][91]+sumram[116][92]+sumram[116][93]+sumram[116][94]+sumram[116][95]+sumram[116][96]+sumram[116][97]+sumram[116][98]+sumram[116][99]+sumram[116][100]+sumram[116][101]+sumram[116][102]+sumram[116][103]+sumram[116][104]+sumram[116][105]+sumram[116][106]+sumram[116][107]+sumram[116][108]+sumram[116][109]+sumram[116][110]+sumram[116][111]+sumram[116][112]+sumram[116][113]+sumram[116][114]+sumram[116][115]+sumram[116][116]+sumram[116][117]+sumram[116][118]+sumram[116][119]+sumram[116][120]+sumram[116][121]+sumram[116][122]+sumram[116][123]+sumram[116][124]+sumram[116][125]+sumram[116][126]+sumram[116][127]+sumram[116][128]+sumram[116][129]+sumram[116][130]+sumram[116][131]+sumram[116][132]+sumram[116][133]+sumram[116][134]+sumram[116][135]+sumram[116][136];
    assign sumcache[117]=sumram[117][0]+sumram[117][1]+sumram[117][2]+sumram[117][3]+sumram[117][4]+sumram[117][5]+sumram[117][6]+sumram[117][7]+sumram[117][8]+sumram[117][9]+sumram[117][10]+sumram[117][11]+sumram[117][12]+sumram[117][13]+sumram[117][14]+sumram[117][15]+sumram[117][16]+sumram[117][17]+sumram[117][18]+sumram[117][19]+sumram[117][20]+sumram[117][21]+sumram[117][22]+sumram[117][23]+sumram[117][24]+sumram[117][25]+sumram[117][26]+sumram[117][27]+sumram[117][28]+sumram[117][29]+sumram[117][30]+sumram[117][31]+sumram[117][32]+sumram[117][33]+sumram[117][34]+sumram[117][35]+sumram[117][36]+sumram[117][37]+sumram[117][38]+sumram[117][39]+sumram[117][40]+sumram[117][41]+sumram[117][42]+sumram[117][43]+sumram[117][44]+sumram[117][45]+sumram[117][46]+sumram[117][47]+sumram[117][48]+sumram[117][49]+sumram[117][50]+sumram[117][51]+sumram[117][52]+sumram[117][53]+sumram[117][54]+sumram[117][55]+sumram[117][56]+sumram[117][57]+sumram[117][58]+sumram[117][59]+sumram[117][60]+sumram[117][61]+sumram[117][62]+sumram[117][63]+sumram[117][64]+sumram[117][65]+sumram[117][66]+sumram[117][67]+sumram[117][68]+sumram[117][69]+sumram[117][70]+sumram[117][71]+sumram[117][72]+sumram[117][73]+sumram[117][74]+sumram[117][75]+sumram[117][76]+sumram[117][77]+sumram[117][78]+sumram[117][79]+sumram[117][80]+sumram[117][81]+sumram[117][82]+sumram[117][83]+sumram[117][84]+sumram[117][85]+sumram[117][86]+sumram[117][87]+sumram[117][88]+sumram[117][89]+sumram[117][90]+sumram[117][91]+sumram[117][92]+sumram[117][93]+sumram[117][94]+sumram[117][95]+sumram[117][96]+sumram[117][97]+sumram[117][98]+sumram[117][99]+sumram[117][100]+sumram[117][101]+sumram[117][102]+sumram[117][103]+sumram[117][104]+sumram[117][105]+sumram[117][106]+sumram[117][107]+sumram[117][108]+sumram[117][109]+sumram[117][110]+sumram[117][111]+sumram[117][112]+sumram[117][113]+sumram[117][114]+sumram[117][115]+sumram[117][116]+sumram[117][117]+sumram[117][118]+sumram[117][119]+sumram[117][120]+sumram[117][121]+sumram[117][122]+sumram[117][123]+sumram[117][124]+sumram[117][125]+sumram[117][126]+sumram[117][127]+sumram[117][128]+sumram[117][129]+sumram[117][130]+sumram[117][131]+sumram[117][132]+sumram[117][133]+sumram[117][134]+sumram[117][135]+sumram[117][136];
    assign sumcache[118]=sumram[118][0]+sumram[118][1]+sumram[118][2]+sumram[118][3]+sumram[118][4]+sumram[118][5]+sumram[118][6]+sumram[118][7]+sumram[118][8]+sumram[118][9]+sumram[118][10]+sumram[118][11]+sumram[118][12]+sumram[118][13]+sumram[118][14]+sumram[118][15]+sumram[118][16]+sumram[118][17]+sumram[118][18]+sumram[118][19]+sumram[118][20]+sumram[118][21]+sumram[118][22]+sumram[118][23]+sumram[118][24]+sumram[118][25]+sumram[118][26]+sumram[118][27]+sumram[118][28]+sumram[118][29]+sumram[118][30]+sumram[118][31]+sumram[118][32]+sumram[118][33]+sumram[118][34]+sumram[118][35]+sumram[118][36]+sumram[118][37]+sumram[118][38]+sumram[118][39]+sumram[118][40]+sumram[118][41]+sumram[118][42]+sumram[118][43]+sumram[118][44]+sumram[118][45]+sumram[118][46]+sumram[118][47]+sumram[118][48]+sumram[118][49]+sumram[118][50]+sumram[118][51]+sumram[118][52]+sumram[118][53]+sumram[118][54]+sumram[118][55]+sumram[118][56]+sumram[118][57]+sumram[118][58]+sumram[118][59]+sumram[118][60]+sumram[118][61]+sumram[118][62]+sumram[118][63]+sumram[118][64]+sumram[118][65]+sumram[118][66]+sumram[118][67]+sumram[118][68]+sumram[118][69]+sumram[118][70]+sumram[118][71]+sumram[118][72]+sumram[118][73]+sumram[118][74]+sumram[118][75]+sumram[118][76]+sumram[118][77]+sumram[118][78]+sumram[118][79]+sumram[118][80]+sumram[118][81]+sumram[118][82]+sumram[118][83]+sumram[118][84]+sumram[118][85]+sumram[118][86]+sumram[118][87]+sumram[118][88]+sumram[118][89]+sumram[118][90]+sumram[118][91]+sumram[118][92]+sumram[118][93]+sumram[118][94]+sumram[118][95]+sumram[118][96]+sumram[118][97]+sumram[118][98]+sumram[118][99]+sumram[118][100]+sumram[118][101]+sumram[118][102]+sumram[118][103]+sumram[118][104]+sumram[118][105]+sumram[118][106]+sumram[118][107]+sumram[118][108]+sumram[118][109]+sumram[118][110]+sumram[118][111]+sumram[118][112]+sumram[118][113]+sumram[118][114]+sumram[118][115]+sumram[118][116]+sumram[118][117]+sumram[118][118]+sumram[118][119]+sumram[118][120]+sumram[118][121]+sumram[118][122]+sumram[118][123]+sumram[118][124]+sumram[118][125]+sumram[118][126]+sumram[118][127]+sumram[118][128]+sumram[118][129]+sumram[118][130]+sumram[118][131]+sumram[118][132]+sumram[118][133]+sumram[118][134]+sumram[118][135]+sumram[118][136];
    assign sumcache[119]=sumram[119][0]+sumram[119][1]+sumram[119][2]+sumram[119][3]+sumram[119][4]+sumram[119][5]+sumram[119][6]+sumram[119][7]+sumram[119][8]+sumram[119][9]+sumram[119][10]+sumram[119][11]+sumram[119][12]+sumram[119][13]+sumram[119][14]+sumram[119][15]+sumram[119][16]+sumram[119][17]+sumram[119][18]+sumram[119][19]+sumram[119][20]+sumram[119][21]+sumram[119][22]+sumram[119][23]+sumram[119][24]+sumram[119][25]+sumram[119][26]+sumram[119][27]+sumram[119][28]+sumram[119][29]+sumram[119][30]+sumram[119][31]+sumram[119][32]+sumram[119][33]+sumram[119][34]+sumram[119][35]+sumram[119][36]+sumram[119][37]+sumram[119][38]+sumram[119][39]+sumram[119][40]+sumram[119][41]+sumram[119][42]+sumram[119][43]+sumram[119][44]+sumram[119][45]+sumram[119][46]+sumram[119][47]+sumram[119][48]+sumram[119][49]+sumram[119][50]+sumram[119][51]+sumram[119][52]+sumram[119][53]+sumram[119][54]+sumram[119][55]+sumram[119][56]+sumram[119][57]+sumram[119][58]+sumram[119][59]+sumram[119][60]+sumram[119][61]+sumram[119][62]+sumram[119][63]+sumram[119][64]+sumram[119][65]+sumram[119][66]+sumram[119][67]+sumram[119][68]+sumram[119][69]+sumram[119][70]+sumram[119][71]+sumram[119][72]+sumram[119][73]+sumram[119][74]+sumram[119][75]+sumram[119][76]+sumram[119][77]+sumram[119][78]+sumram[119][79]+sumram[119][80]+sumram[119][81]+sumram[119][82]+sumram[119][83]+sumram[119][84]+sumram[119][85]+sumram[119][86]+sumram[119][87]+sumram[119][88]+sumram[119][89]+sumram[119][90]+sumram[119][91]+sumram[119][92]+sumram[119][93]+sumram[119][94]+sumram[119][95]+sumram[119][96]+sumram[119][97]+sumram[119][98]+sumram[119][99]+sumram[119][100]+sumram[119][101]+sumram[119][102]+sumram[119][103]+sumram[119][104]+sumram[119][105]+sumram[119][106]+sumram[119][107]+sumram[119][108]+sumram[119][109]+sumram[119][110]+sumram[119][111]+sumram[119][112]+sumram[119][113]+sumram[119][114]+sumram[119][115]+sumram[119][116]+sumram[119][117]+sumram[119][118]+sumram[119][119]+sumram[119][120]+sumram[119][121]+sumram[119][122]+sumram[119][123]+sumram[119][124]+sumram[119][125]+sumram[119][126]+sumram[119][127]+sumram[119][128]+sumram[119][129]+sumram[119][130]+sumram[119][131]+sumram[119][132]+sumram[119][133]+sumram[119][134]+sumram[119][135]+sumram[119][136];
    assign sumcache[120]=sumram[120][0]+sumram[120][1]+sumram[120][2]+sumram[120][3]+sumram[120][4]+sumram[120][5]+sumram[120][6]+sumram[120][7]+sumram[120][8]+sumram[120][9]+sumram[120][10]+sumram[120][11]+sumram[120][12]+sumram[120][13]+sumram[120][14]+sumram[120][15]+sumram[120][16]+sumram[120][17]+sumram[120][18]+sumram[120][19]+sumram[120][20]+sumram[120][21]+sumram[120][22]+sumram[120][23]+sumram[120][24]+sumram[120][25]+sumram[120][26]+sumram[120][27]+sumram[120][28]+sumram[120][29]+sumram[120][30]+sumram[120][31]+sumram[120][32]+sumram[120][33]+sumram[120][34]+sumram[120][35]+sumram[120][36]+sumram[120][37]+sumram[120][38]+sumram[120][39]+sumram[120][40]+sumram[120][41]+sumram[120][42]+sumram[120][43]+sumram[120][44]+sumram[120][45]+sumram[120][46]+sumram[120][47]+sumram[120][48]+sumram[120][49]+sumram[120][50]+sumram[120][51]+sumram[120][52]+sumram[120][53]+sumram[120][54]+sumram[120][55]+sumram[120][56]+sumram[120][57]+sumram[120][58]+sumram[120][59]+sumram[120][60]+sumram[120][61]+sumram[120][62]+sumram[120][63]+sumram[120][64]+sumram[120][65]+sumram[120][66]+sumram[120][67]+sumram[120][68]+sumram[120][69]+sumram[120][70]+sumram[120][71]+sumram[120][72]+sumram[120][73]+sumram[120][74]+sumram[120][75]+sumram[120][76]+sumram[120][77]+sumram[120][78]+sumram[120][79]+sumram[120][80]+sumram[120][81]+sumram[120][82]+sumram[120][83]+sumram[120][84]+sumram[120][85]+sumram[120][86]+sumram[120][87]+sumram[120][88]+sumram[120][89]+sumram[120][90]+sumram[120][91]+sumram[120][92]+sumram[120][93]+sumram[120][94]+sumram[120][95]+sumram[120][96]+sumram[120][97]+sumram[120][98]+sumram[120][99]+sumram[120][100]+sumram[120][101]+sumram[120][102]+sumram[120][103]+sumram[120][104]+sumram[120][105]+sumram[120][106]+sumram[120][107]+sumram[120][108]+sumram[120][109]+sumram[120][110]+sumram[120][111]+sumram[120][112]+sumram[120][113]+sumram[120][114]+sumram[120][115]+sumram[120][116]+sumram[120][117]+sumram[120][118]+sumram[120][119]+sumram[120][120]+sumram[120][121]+sumram[120][122]+sumram[120][123]+sumram[120][124]+sumram[120][125]+sumram[120][126]+sumram[120][127]+sumram[120][128]+sumram[120][129]+sumram[120][130]+sumram[120][131]+sumram[120][132]+sumram[120][133]+sumram[120][134]+sumram[120][135]+sumram[120][136];
    assign sumcache[121]=sumram[121][0]+sumram[121][1]+sumram[121][2]+sumram[121][3]+sumram[121][4]+sumram[121][5]+sumram[121][6]+sumram[121][7]+sumram[121][8]+sumram[121][9]+sumram[121][10]+sumram[121][11]+sumram[121][12]+sumram[121][13]+sumram[121][14]+sumram[121][15]+sumram[121][16]+sumram[121][17]+sumram[121][18]+sumram[121][19]+sumram[121][20]+sumram[121][21]+sumram[121][22]+sumram[121][23]+sumram[121][24]+sumram[121][25]+sumram[121][26]+sumram[121][27]+sumram[121][28]+sumram[121][29]+sumram[121][30]+sumram[121][31]+sumram[121][32]+sumram[121][33]+sumram[121][34]+sumram[121][35]+sumram[121][36]+sumram[121][37]+sumram[121][38]+sumram[121][39]+sumram[121][40]+sumram[121][41]+sumram[121][42]+sumram[121][43]+sumram[121][44]+sumram[121][45]+sumram[121][46]+sumram[121][47]+sumram[121][48]+sumram[121][49]+sumram[121][50]+sumram[121][51]+sumram[121][52]+sumram[121][53]+sumram[121][54]+sumram[121][55]+sumram[121][56]+sumram[121][57]+sumram[121][58]+sumram[121][59]+sumram[121][60]+sumram[121][61]+sumram[121][62]+sumram[121][63]+sumram[121][64]+sumram[121][65]+sumram[121][66]+sumram[121][67]+sumram[121][68]+sumram[121][69]+sumram[121][70]+sumram[121][71]+sumram[121][72]+sumram[121][73]+sumram[121][74]+sumram[121][75]+sumram[121][76]+sumram[121][77]+sumram[121][78]+sumram[121][79]+sumram[121][80]+sumram[121][81]+sumram[121][82]+sumram[121][83]+sumram[121][84]+sumram[121][85]+sumram[121][86]+sumram[121][87]+sumram[121][88]+sumram[121][89]+sumram[121][90]+sumram[121][91]+sumram[121][92]+sumram[121][93]+sumram[121][94]+sumram[121][95]+sumram[121][96]+sumram[121][97]+sumram[121][98]+sumram[121][99]+sumram[121][100]+sumram[121][101]+sumram[121][102]+sumram[121][103]+sumram[121][104]+sumram[121][105]+sumram[121][106]+sumram[121][107]+sumram[121][108]+sumram[121][109]+sumram[121][110]+sumram[121][111]+sumram[121][112]+sumram[121][113]+sumram[121][114]+sumram[121][115]+sumram[121][116]+sumram[121][117]+sumram[121][118]+sumram[121][119]+sumram[121][120]+sumram[121][121]+sumram[121][122]+sumram[121][123]+sumram[121][124]+sumram[121][125]+sumram[121][126]+sumram[121][127]+sumram[121][128]+sumram[121][129]+sumram[121][130]+sumram[121][131]+sumram[121][132]+sumram[121][133]+sumram[121][134]+sumram[121][135]+sumram[121][136];
    assign sumcache[122]=sumram[122][0]+sumram[122][1]+sumram[122][2]+sumram[122][3]+sumram[122][4]+sumram[122][5]+sumram[122][6]+sumram[122][7]+sumram[122][8]+sumram[122][9]+sumram[122][10]+sumram[122][11]+sumram[122][12]+sumram[122][13]+sumram[122][14]+sumram[122][15]+sumram[122][16]+sumram[122][17]+sumram[122][18]+sumram[122][19]+sumram[122][20]+sumram[122][21]+sumram[122][22]+sumram[122][23]+sumram[122][24]+sumram[122][25]+sumram[122][26]+sumram[122][27]+sumram[122][28]+sumram[122][29]+sumram[122][30]+sumram[122][31]+sumram[122][32]+sumram[122][33]+sumram[122][34]+sumram[122][35]+sumram[122][36]+sumram[122][37]+sumram[122][38]+sumram[122][39]+sumram[122][40]+sumram[122][41]+sumram[122][42]+sumram[122][43]+sumram[122][44]+sumram[122][45]+sumram[122][46]+sumram[122][47]+sumram[122][48]+sumram[122][49]+sumram[122][50]+sumram[122][51]+sumram[122][52]+sumram[122][53]+sumram[122][54]+sumram[122][55]+sumram[122][56]+sumram[122][57]+sumram[122][58]+sumram[122][59]+sumram[122][60]+sumram[122][61]+sumram[122][62]+sumram[122][63]+sumram[122][64]+sumram[122][65]+sumram[122][66]+sumram[122][67]+sumram[122][68]+sumram[122][69]+sumram[122][70]+sumram[122][71]+sumram[122][72]+sumram[122][73]+sumram[122][74]+sumram[122][75]+sumram[122][76]+sumram[122][77]+sumram[122][78]+sumram[122][79]+sumram[122][80]+sumram[122][81]+sumram[122][82]+sumram[122][83]+sumram[122][84]+sumram[122][85]+sumram[122][86]+sumram[122][87]+sumram[122][88]+sumram[122][89]+sumram[122][90]+sumram[122][91]+sumram[122][92]+sumram[122][93]+sumram[122][94]+sumram[122][95]+sumram[122][96]+sumram[122][97]+sumram[122][98]+sumram[122][99]+sumram[122][100]+sumram[122][101]+sumram[122][102]+sumram[122][103]+sumram[122][104]+sumram[122][105]+sumram[122][106]+sumram[122][107]+sumram[122][108]+sumram[122][109]+sumram[122][110]+sumram[122][111]+sumram[122][112]+sumram[122][113]+sumram[122][114]+sumram[122][115]+sumram[122][116]+sumram[122][117]+sumram[122][118]+sumram[122][119]+sumram[122][120]+sumram[122][121]+sumram[122][122]+sumram[122][123]+sumram[122][124]+sumram[122][125]+sumram[122][126]+sumram[122][127]+sumram[122][128]+sumram[122][129]+sumram[122][130]+sumram[122][131]+sumram[122][132]+sumram[122][133]+sumram[122][134]+sumram[122][135]+sumram[122][136];
    assign sumcache[123]=sumram[123][0]+sumram[123][1]+sumram[123][2]+sumram[123][3]+sumram[123][4]+sumram[123][5]+sumram[123][6]+sumram[123][7]+sumram[123][8]+sumram[123][9]+sumram[123][10]+sumram[123][11]+sumram[123][12]+sumram[123][13]+sumram[123][14]+sumram[123][15]+sumram[123][16]+sumram[123][17]+sumram[123][18]+sumram[123][19]+sumram[123][20]+sumram[123][21]+sumram[123][22]+sumram[123][23]+sumram[123][24]+sumram[123][25]+sumram[123][26]+sumram[123][27]+sumram[123][28]+sumram[123][29]+sumram[123][30]+sumram[123][31]+sumram[123][32]+sumram[123][33]+sumram[123][34]+sumram[123][35]+sumram[123][36]+sumram[123][37]+sumram[123][38]+sumram[123][39]+sumram[123][40]+sumram[123][41]+sumram[123][42]+sumram[123][43]+sumram[123][44]+sumram[123][45]+sumram[123][46]+sumram[123][47]+sumram[123][48]+sumram[123][49]+sumram[123][50]+sumram[123][51]+sumram[123][52]+sumram[123][53]+sumram[123][54]+sumram[123][55]+sumram[123][56]+sumram[123][57]+sumram[123][58]+sumram[123][59]+sumram[123][60]+sumram[123][61]+sumram[123][62]+sumram[123][63]+sumram[123][64]+sumram[123][65]+sumram[123][66]+sumram[123][67]+sumram[123][68]+sumram[123][69]+sumram[123][70]+sumram[123][71]+sumram[123][72]+sumram[123][73]+sumram[123][74]+sumram[123][75]+sumram[123][76]+sumram[123][77]+sumram[123][78]+sumram[123][79]+sumram[123][80]+sumram[123][81]+sumram[123][82]+sumram[123][83]+sumram[123][84]+sumram[123][85]+sumram[123][86]+sumram[123][87]+sumram[123][88]+sumram[123][89]+sumram[123][90]+sumram[123][91]+sumram[123][92]+sumram[123][93]+sumram[123][94]+sumram[123][95]+sumram[123][96]+sumram[123][97]+sumram[123][98]+sumram[123][99]+sumram[123][100]+sumram[123][101]+sumram[123][102]+sumram[123][103]+sumram[123][104]+sumram[123][105]+sumram[123][106]+sumram[123][107]+sumram[123][108]+sumram[123][109]+sumram[123][110]+sumram[123][111]+sumram[123][112]+sumram[123][113]+sumram[123][114]+sumram[123][115]+sumram[123][116]+sumram[123][117]+sumram[123][118]+sumram[123][119]+sumram[123][120]+sumram[123][121]+sumram[123][122]+sumram[123][123]+sumram[123][124]+sumram[123][125]+sumram[123][126]+sumram[123][127]+sumram[123][128]+sumram[123][129]+sumram[123][130]+sumram[123][131]+sumram[123][132]+sumram[123][133]+sumram[123][134]+sumram[123][135]+sumram[123][136];
    assign sumcache[124]=sumram[124][0]+sumram[124][1]+sumram[124][2]+sumram[124][3]+sumram[124][4]+sumram[124][5]+sumram[124][6]+sumram[124][7]+sumram[124][8]+sumram[124][9]+sumram[124][10]+sumram[124][11]+sumram[124][12]+sumram[124][13]+sumram[124][14]+sumram[124][15]+sumram[124][16]+sumram[124][17]+sumram[124][18]+sumram[124][19]+sumram[124][20]+sumram[124][21]+sumram[124][22]+sumram[124][23]+sumram[124][24]+sumram[124][25]+sumram[124][26]+sumram[124][27]+sumram[124][28]+sumram[124][29]+sumram[124][30]+sumram[124][31]+sumram[124][32]+sumram[124][33]+sumram[124][34]+sumram[124][35]+sumram[124][36]+sumram[124][37]+sumram[124][38]+sumram[124][39]+sumram[124][40]+sumram[124][41]+sumram[124][42]+sumram[124][43]+sumram[124][44]+sumram[124][45]+sumram[124][46]+sumram[124][47]+sumram[124][48]+sumram[124][49]+sumram[124][50]+sumram[124][51]+sumram[124][52]+sumram[124][53]+sumram[124][54]+sumram[124][55]+sumram[124][56]+sumram[124][57]+sumram[124][58]+sumram[124][59]+sumram[124][60]+sumram[124][61]+sumram[124][62]+sumram[124][63]+sumram[124][64]+sumram[124][65]+sumram[124][66]+sumram[124][67]+sumram[124][68]+sumram[124][69]+sumram[124][70]+sumram[124][71]+sumram[124][72]+sumram[124][73]+sumram[124][74]+sumram[124][75]+sumram[124][76]+sumram[124][77]+sumram[124][78]+sumram[124][79]+sumram[124][80]+sumram[124][81]+sumram[124][82]+sumram[124][83]+sumram[124][84]+sumram[124][85]+sumram[124][86]+sumram[124][87]+sumram[124][88]+sumram[124][89]+sumram[124][90]+sumram[124][91]+sumram[124][92]+sumram[124][93]+sumram[124][94]+sumram[124][95]+sumram[124][96]+sumram[124][97]+sumram[124][98]+sumram[124][99]+sumram[124][100]+sumram[124][101]+sumram[124][102]+sumram[124][103]+sumram[124][104]+sumram[124][105]+sumram[124][106]+sumram[124][107]+sumram[124][108]+sumram[124][109]+sumram[124][110]+sumram[124][111]+sumram[124][112]+sumram[124][113]+sumram[124][114]+sumram[124][115]+sumram[124][116]+sumram[124][117]+sumram[124][118]+sumram[124][119]+sumram[124][120]+sumram[124][121]+sumram[124][122]+sumram[124][123]+sumram[124][124]+sumram[124][125]+sumram[124][126]+sumram[124][127]+sumram[124][128]+sumram[124][129]+sumram[124][130]+sumram[124][131]+sumram[124][132]+sumram[124][133]+sumram[124][134]+sumram[124][135]+sumram[124][136];
    assign sumcache[125]=sumram[125][0]+sumram[125][1]+sumram[125][2]+sumram[125][3]+sumram[125][4]+sumram[125][5]+sumram[125][6]+sumram[125][7]+sumram[125][8]+sumram[125][9]+sumram[125][10]+sumram[125][11]+sumram[125][12]+sumram[125][13]+sumram[125][14]+sumram[125][15]+sumram[125][16]+sumram[125][17]+sumram[125][18]+sumram[125][19]+sumram[125][20]+sumram[125][21]+sumram[125][22]+sumram[125][23]+sumram[125][24]+sumram[125][25]+sumram[125][26]+sumram[125][27]+sumram[125][28]+sumram[125][29]+sumram[125][30]+sumram[125][31]+sumram[125][32]+sumram[125][33]+sumram[125][34]+sumram[125][35]+sumram[125][36]+sumram[125][37]+sumram[125][38]+sumram[125][39]+sumram[125][40]+sumram[125][41]+sumram[125][42]+sumram[125][43]+sumram[125][44]+sumram[125][45]+sumram[125][46]+sumram[125][47]+sumram[125][48]+sumram[125][49]+sumram[125][50]+sumram[125][51]+sumram[125][52]+sumram[125][53]+sumram[125][54]+sumram[125][55]+sumram[125][56]+sumram[125][57]+sumram[125][58]+sumram[125][59]+sumram[125][60]+sumram[125][61]+sumram[125][62]+sumram[125][63]+sumram[125][64]+sumram[125][65]+sumram[125][66]+sumram[125][67]+sumram[125][68]+sumram[125][69]+sumram[125][70]+sumram[125][71]+sumram[125][72]+sumram[125][73]+sumram[125][74]+sumram[125][75]+sumram[125][76]+sumram[125][77]+sumram[125][78]+sumram[125][79]+sumram[125][80]+sumram[125][81]+sumram[125][82]+sumram[125][83]+sumram[125][84]+sumram[125][85]+sumram[125][86]+sumram[125][87]+sumram[125][88]+sumram[125][89]+sumram[125][90]+sumram[125][91]+sumram[125][92]+sumram[125][93]+sumram[125][94]+sumram[125][95]+sumram[125][96]+sumram[125][97]+sumram[125][98]+sumram[125][99]+sumram[125][100]+sumram[125][101]+sumram[125][102]+sumram[125][103]+sumram[125][104]+sumram[125][105]+sumram[125][106]+sumram[125][107]+sumram[125][108]+sumram[125][109]+sumram[125][110]+sumram[125][111]+sumram[125][112]+sumram[125][113]+sumram[125][114]+sumram[125][115]+sumram[125][116]+sumram[125][117]+sumram[125][118]+sumram[125][119]+sumram[125][120]+sumram[125][121]+sumram[125][122]+sumram[125][123]+sumram[125][124]+sumram[125][125]+sumram[125][126]+sumram[125][127]+sumram[125][128]+sumram[125][129]+sumram[125][130]+sumram[125][131]+sumram[125][132]+sumram[125][133]+sumram[125][134]+sumram[125][135]+sumram[125][136];
    assign sumcache[126]=sumram[126][0]+sumram[126][1]+sumram[126][2]+sumram[126][3]+sumram[126][4]+sumram[126][5]+sumram[126][6]+sumram[126][7]+sumram[126][8]+sumram[126][9]+sumram[126][10]+sumram[126][11]+sumram[126][12]+sumram[126][13]+sumram[126][14]+sumram[126][15]+sumram[126][16]+sumram[126][17]+sumram[126][18]+sumram[126][19]+sumram[126][20]+sumram[126][21]+sumram[126][22]+sumram[126][23]+sumram[126][24]+sumram[126][25]+sumram[126][26]+sumram[126][27]+sumram[126][28]+sumram[126][29]+sumram[126][30]+sumram[126][31]+sumram[126][32]+sumram[126][33]+sumram[126][34]+sumram[126][35]+sumram[126][36]+sumram[126][37]+sumram[126][38]+sumram[126][39]+sumram[126][40]+sumram[126][41]+sumram[126][42]+sumram[126][43]+sumram[126][44]+sumram[126][45]+sumram[126][46]+sumram[126][47]+sumram[126][48]+sumram[126][49]+sumram[126][50]+sumram[126][51]+sumram[126][52]+sumram[126][53]+sumram[126][54]+sumram[126][55]+sumram[126][56]+sumram[126][57]+sumram[126][58]+sumram[126][59]+sumram[126][60]+sumram[126][61]+sumram[126][62]+sumram[126][63]+sumram[126][64]+sumram[126][65]+sumram[126][66]+sumram[126][67]+sumram[126][68]+sumram[126][69]+sumram[126][70]+sumram[126][71]+sumram[126][72]+sumram[126][73]+sumram[126][74]+sumram[126][75]+sumram[126][76]+sumram[126][77]+sumram[126][78]+sumram[126][79]+sumram[126][80]+sumram[126][81]+sumram[126][82]+sumram[126][83]+sumram[126][84]+sumram[126][85]+sumram[126][86]+sumram[126][87]+sumram[126][88]+sumram[126][89]+sumram[126][90]+sumram[126][91]+sumram[126][92]+sumram[126][93]+sumram[126][94]+sumram[126][95]+sumram[126][96]+sumram[126][97]+sumram[126][98]+sumram[126][99]+sumram[126][100]+sumram[126][101]+sumram[126][102]+sumram[126][103]+sumram[126][104]+sumram[126][105]+sumram[126][106]+sumram[126][107]+sumram[126][108]+sumram[126][109]+sumram[126][110]+sumram[126][111]+sumram[126][112]+sumram[126][113]+sumram[126][114]+sumram[126][115]+sumram[126][116]+sumram[126][117]+sumram[126][118]+sumram[126][119]+sumram[126][120]+sumram[126][121]+sumram[126][122]+sumram[126][123]+sumram[126][124]+sumram[126][125]+sumram[126][126]+sumram[126][127]+sumram[126][128]+sumram[126][129]+sumram[126][130]+sumram[126][131]+sumram[126][132]+sumram[126][133]+sumram[126][134]+sumram[126][135]+sumram[126][136];
    assign sumcache[127]=sumram[127][0]+sumram[127][1]+sumram[127][2]+sumram[127][3]+sumram[127][4]+sumram[127][5]+sumram[127][6]+sumram[127][7]+sumram[127][8]+sumram[127][9]+sumram[127][10]+sumram[127][11]+sumram[127][12]+sumram[127][13]+sumram[127][14]+sumram[127][15]+sumram[127][16]+sumram[127][17]+sumram[127][18]+sumram[127][19]+sumram[127][20]+sumram[127][21]+sumram[127][22]+sumram[127][23]+sumram[127][24]+sumram[127][25]+sumram[127][26]+sumram[127][27]+sumram[127][28]+sumram[127][29]+sumram[127][30]+sumram[127][31]+sumram[127][32]+sumram[127][33]+sumram[127][34]+sumram[127][35]+sumram[127][36]+sumram[127][37]+sumram[127][38]+sumram[127][39]+sumram[127][40]+sumram[127][41]+sumram[127][42]+sumram[127][43]+sumram[127][44]+sumram[127][45]+sumram[127][46]+sumram[127][47]+sumram[127][48]+sumram[127][49]+sumram[127][50]+sumram[127][51]+sumram[127][52]+sumram[127][53]+sumram[127][54]+sumram[127][55]+sumram[127][56]+sumram[127][57]+sumram[127][58]+sumram[127][59]+sumram[127][60]+sumram[127][61]+sumram[127][62]+sumram[127][63]+sumram[127][64]+sumram[127][65]+sumram[127][66]+sumram[127][67]+sumram[127][68]+sumram[127][69]+sumram[127][70]+sumram[127][71]+sumram[127][72]+sumram[127][73]+sumram[127][74]+sumram[127][75]+sumram[127][76]+sumram[127][77]+sumram[127][78]+sumram[127][79]+sumram[127][80]+sumram[127][81]+sumram[127][82]+sumram[127][83]+sumram[127][84]+sumram[127][85]+sumram[127][86]+sumram[127][87]+sumram[127][88]+sumram[127][89]+sumram[127][90]+sumram[127][91]+sumram[127][92]+sumram[127][93]+sumram[127][94]+sumram[127][95]+sumram[127][96]+sumram[127][97]+sumram[127][98]+sumram[127][99]+sumram[127][100]+sumram[127][101]+sumram[127][102]+sumram[127][103]+sumram[127][104]+sumram[127][105]+sumram[127][106]+sumram[127][107]+sumram[127][108]+sumram[127][109]+sumram[127][110]+sumram[127][111]+sumram[127][112]+sumram[127][113]+sumram[127][114]+sumram[127][115]+sumram[127][116]+sumram[127][117]+sumram[127][118]+sumram[127][119]+sumram[127][120]+sumram[127][121]+sumram[127][122]+sumram[127][123]+sumram[127][124]+sumram[127][125]+sumram[127][126]+sumram[127][127]+sumram[127][128]+sumram[127][129]+sumram[127][130]+sumram[127][131]+sumram[127][132]+sumram[127][133]+sumram[127][134]+sumram[127][135]+sumram[127][136];
    assign sumcache[128]=sumram[128][0]+sumram[128][1]+sumram[128][2]+sumram[128][3]+sumram[128][4]+sumram[128][5]+sumram[128][6]+sumram[128][7]+sumram[128][8]+sumram[128][9]+sumram[128][10]+sumram[128][11]+sumram[128][12]+sumram[128][13]+sumram[128][14]+sumram[128][15]+sumram[128][16]+sumram[128][17]+sumram[128][18]+sumram[128][19]+sumram[128][20]+sumram[128][21]+sumram[128][22]+sumram[128][23]+sumram[128][24]+sumram[128][25]+sumram[128][26]+sumram[128][27]+sumram[128][28]+sumram[128][29]+sumram[128][30]+sumram[128][31]+sumram[128][32]+sumram[128][33]+sumram[128][34]+sumram[128][35]+sumram[128][36]+sumram[128][37]+sumram[128][38]+sumram[128][39]+sumram[128][40]+sumram[128][41]+sumram[128][42]+sumram[128][43]+sumram[128][44]+sumram[128][45]+sumram[128][46]+sumram[128][47]+sumram[128][48]+sumram[128][49]+sumram[128][50]+sumram[128][51]+sumram[128][52]+sumram[128][53]+sumram[128][54]+sumram[128][55]+sumram[128][56]+sumram[128][57]+sumram[128][58]+sumram[128][59]+sumram[128][60]+sumram[128][61]+sumram[128][62]+sumram[128][63]+sumram[128][64]+sumram[128][65]+sumram[128][66]+sumram[128][67]+sumram[128][68]+sumram[128][69]+sumram[128][70]+sumram[128][71]+sumram[128][72]+sumram[128][73]+sumram[128][74]+sumram[128][75]+sumram[128][76]+sumram[128][77]+sumram[128][78]+sumram[128][79]+sumram[128][80]+sumram[128][81]+sumram[128][82]+sumram[128][83]+sumram[128][84]+sumram[128][85]+sumram[128][86]+sumram[128][87]+sumram[128][88]+sumram[128][89]+sumram[128][90]+sumram[128][91]+sumram[128][92]+sumram[128][93]+sumram[128][94]+sumram[128][95]+sumram[128][96]+sumram[128][97]+sumram[128][98]+sumram[128][99]+sumram[128][100]+sumram[128][101]+sumram[128][102]+sumram[128][103]+sumram[128][104]+sumram[128][105]+sumram[128][106]+sumram[128][107]+sumram[128][108]+sumram[128][109]+sumram[128][110]+sumram[128][111]+sumram[128][112]+sumram[128][113]+sumram[128][114]+sumram[128][115]+sumram[128][116]+sumram[128][117]+sumram[128][118]+sumram[128][119]+sumram[128][120]+sumram[128][121]+sumram[128][122]+sumram[128][123]+sumram[128][124]+sumram[128][125]+sumram[128][126]+sumram[128][127]+sumram[128][128]+sumram[128][129]+sumram[128][130]+sumram[128][131]+sumram[128][132]+sumram[128][133]+sumram[128][134]+sumram[128][135]+sumram[128][136];
    assign sumcache[129]=sumram[129][0]+sumram[129][1]+sumram[129][2]+sumram[129][3]+sumram[129][4]+sumram[129][5]+sumram[129][6]+sumram[129][7]+sumram[129][8]+sumram[129][9]+sumram[129][10]+sumram[129][11]+sumram[129][12]+sumram[129][13]+sumram[129][14]+sumram[129][15]+sumram[129][16]+sumram[129][17]+sumram[129][18]+sumram[129][19]+sumram[129][20]+sumram[129][21]+sumram[129][22]+sumram[129][23]+sumram[129][24]+sumram[129][25]+sumram[129][26]+sumram[129][27]+sumram[129][28]+sumram[129][29]+sumram[129][30]+sumram[129][31]+sumram[129][32]+sumram[129][33]+sumram[129][34]+sumram[129][35]+sumram[129][36]+sumram[129][37]+sumram[129][38]+sumram[129][39]+sumram[129][40]+sumram[129][41]+sumram[129][42]+sumram[129][43]+sumram[129][44]+sumram[129][45]+sumram[129][46]+sumram[129][47]+sumram[129][48]+sumram[129][49]+sumram[129][50]+sumram[129][51]+sumram[129][52]+sumram[129][53]+sumram[129][54]+sumram[129][55]+sumram[129][56]+sumram[129][57]+sumram[129][58]+sumram[129][59]+sumram[129][60]+sumram[129][61]+sumram[129][62]+sumram[129][63]+sumram[129][64]+sumram[129][65]+sumram[129][66]+sumram[129][67]+sumram[129][68]+sumram[129][69]+sumram[129][70]+sumram[129][71]+sumram[129][72]+sumram[129][73]+sumram[129][74]+sumram[129][75]+sumram[129][76]+sumram[129][77]+sumram[129][78]+sumram[129][79]+sumram[129][80]+sumram[129][81]+sumram[129][82]+sumram[129][83]+sumram[129][84]+sumram[129][85]+sumram[129][86]+sumram[129][87]+sumram[129][88]+sumram[129][89]+sumram[129][90]+sumram[129][91]+sumram[129][92]+sumram[129][93]+sumram[129][94]+sumram[129][95]+sumram[129][96]+sumram[129][97]+sumram[129][98]+sumram[129][99]+sumram[129][100]+sumram[129][101]+sumram[129][102]+sumram[129][103]+sumram[129][104]+sumram[129][105]+sumram[129][106]+sumram[129][107]+sumram[129][108]+sumram[129][109]+sumram[129][110]+sumram[129][111]+sumram[129][112]+sumram[129][113]+sumram[129][114]+sumram[129][115]+sumram[129][116]+sumram[129][117]+sumram[129][118]+sumram[129][119]+sumram[129][120]+sumram[129][121]+sumram[129][122]+sumram[129][123]+sumram[129][124]+sumram[129][125]+sumram[129][126]+sumram[129][127]+sumram[129][128]+sumram[129][129]+sumram[129][130]+sumram[129][131]+sumram[129][132]+sumram[129][133]+sumram[129][134]+sumram[129][135]+sumram[129][136];
    assign sumcache[130]=sumram[130][0]+sumram[130][1]+sumram[130][2]+sumram[130][3]+sumram[130][4]+sumram[130][5]+sumram[130][6]+sumram[130][7]+sumram[130][8]+sumram[130][9]+sumram[130][10]+sumram[130][11]+sumram[130][12]+sumram[130][13]+sumram[130][14]+sumram[130][15]+sumram[130][16]+sumram[130][17]+sumram[130][18]+sumram[130][19]+sumram[130][20]+sumram[130][21]+sumram[130][22]+sumram[130][23]+sumram[130][24]+sumram[130][25]+sumram[130][26]+sumram[130][27]+sumram[130][28]+sumram[130][29]+sumram[130][30]+sumram[130][31]+sumram[130][32]+sumram[130][33]+sumram[130][34]+sumram[130][35]+sumram[130][36]+sumram[130][37]+sumram[130][38]+sumram[130][39]+sumram[130][40]+sumram[130][41]+sumram[130][42]+sumram[130][43]+sumram[130][44]+sumram[130][45]+sumram[130][46]+sumram[130][47]+sumram[130][48]+sumram[130][49]+sumram[130][50]+sumram[130][51]+sumram[130][52]+sumram[130][53]+sumram[130][54]+sumram[130][55]+sumram[130][56]+sumram[130][57]+sumram[130][58]+sumram[130][59]+sumram[130][60]+sumram[130][61]+sumram[130][62]+sumram[130][63]+sumram[130][64]+sumram[130][65]+sumram[130][66]+sumram[130][67]+sumram[130][68]+sumram[130][69]+sumram[130][70]+sumram[130][71]+sumram[130][72]+sumram[130][73]+sumram[130][74]+sumram[130][75]+sumram[130][76]+sumram[130][77]+sumram[130][78]+sumram[130][79]+sumram[130][80]+sumram[130][81]+sumram[130][82]+sumram[130][83]+sumram[130][84]+sumram[130][85]+sumram[130][86]+sumram[130][87]+sumram[130][88]+sumram[130][89]+sumram[130][90]+sumram[130][91]+sumram[130][92]+sumram[130][93]+sumram[130][94]+sumram[130][95]+sumram[130][96]+sumram[130][97]+sumram[130][98]+sumram[130][99]+sumram[130][100]+sumram[130][101]+sumram[130][102]+sumram[130][103]+sumram[130][104]+sumram[130][105]+sumram[130][106]+sumram[130][107]+sumram[130][108]+sumram[130][109]+sumram[130][110]+sumram[130][111]+sumram[130][112]+sumram[130][113]+sumram[130][114]+sumram[130][115]+sumram[130][116]+sumram[130][117]+sumram[130][118]+sumram[130][119]+sumram[130][120]+sumram[130][121]+sumram[130][122]+sumram[130][123]+sumram[130][124]+sumram[130][125]+sumram[130][126]+sumram[130][127]+sumram[130][128]+sumram[130][129]+sumram[130][130]+sumram[130][131]+sumram[130][132]+sumram[130][133]+sumram[130][134]+sumram[130][135]+sumram[130][136];
    assign sumcache[131]=sumram[131][0]+sumram[131][1]+sumram[131][2]+sumram[131][3]+sumram[131][4]+sumram[131][5]+sumram[131][6]+sumram[131][7]+sumram[131][8]+sumram[131][9]+sumram[131][10]+sumram[131][11]+sumram[131][12]+sumram[131][13]+sumram[131][14]+sumram[131][15]+sumram[131][16]+sumram[131][17]+sumram[131][18]+sumram[131][19]+sumram[131][20]+sumram[131][21]+sumram[131][22]+sumram[131][23]+sumram[131][24]+sumram[131][25]+sumram[131][26]+sumram[131][27]+sumram[131][28]+sumram[131][29]+sumram[131][30]+sumram[131][31]+sumram[131][32]+sumram[131][33]+sumram[131][34]+sumram[131][35]+sumram[131][36]+sumram[131][37]+sumram[131][38]+sumram[131][39]+sumram[131][40]+sumram[131][41]+sumram[131][42]+sumram[131][43]+sumram[131][44]+sumram[131][45]+sumram[131][46]+sumram[131][47]+sumram[131][48]+sumram[131][49]+sumram[131][50]+sumram[131][51]+sumram[131][52]+sumram[131][53]+sumram[131][54]+sumram[131][55]+sumram[131][56]+sumram[131][57]+sumram[131][58]+sumram[131][59]+sumram[131][60]+sumram[131][61]+sumram[131][62]+sumram[131][63]+sumram[131][64]+sumram[131][65]+sumram[131][66]+sumram[131][67]+sumram[131][68]+sumram[131][69]+sumram[131][70]+sumram[131][71]+sumram[131][72]+sumram[131][73]+sumram[131][74]+sumram[131][75]+sumram[131][76]+sumram[131][77]+sumram[131][78]+sumram[131][79]+sumram[131][80]+sumram[131][81]+sumram[131][82]+sumram[131][83]+sumram[131][84]+sumram[131][85]+sumram[131][86]+sumram[131][87]+sumram[131][88]+sumram[131][89]+sumram[131][90]+sumram[131][91]+sumram[131][92]+sumram[131][93]+sumram[131][94]+sumram[131][95]+sumram[131][96]+sumram[131][97]+sumram[131][98]+sumram[131][99]+sumram[131][100]+sumram[131][101]+sumram[131][102]+sumram[131][103]+sumram[131][104]+sumram[131][105]+sumram[131][106]+sumram[131][107]+sumram[131][108]+sumram[131][109]+sumram[131][110]+sumram[131][111]+sumram[131][112]+sumram[131][113]+sumram[131][114]+sumram[131][115]+sumram[131][116]+sumram[131][117]+sumram[131][118]+sumram[131][119]+sumram[131][120]+sumram[131][121]+sumram[131][122]+sumram[131][123]+sumram[131][124]+sumram[131][125]+sumram[131][126]+sumram[131][127]+sumram[131][128]+sumram[131][129]+sumram[131][130]+sumram[131][131]+sumram[131][132]+sumram[131][133]+sumram[131][134]+sumram[131][135]+sumram[131][136];
    assign sumcache[132]=sumram[132][0]+sumram[132][1]+sumram[132][2]+sumram[132][3]+sumram[132][4]+sumram[132][5]+sumram[132][6]+sumram[132][7]+sumram[132][8]+sumram[132][9]+sumram[132][10]+sumram[132][11]+sumram[132][12]+sumram[132][13]+sumram[132][14]+sumram[132][15]+sumram[132][16]+sumram[132][17]+sumram[132][18]+sumram[132][19]+sumram[132][20]+sumram[132][21]+sumram[132][22]+sumram[132][23]+sumram[132][24]+sumram[132][25]+sumram[132][26]+sumram[132][27]+sumram[132][28]+sumram[132][29]+sumram[132][30]+sumram[132][31]+sumram[132][32]+sumram[132][33]+sumram[132][34]+sumram[132][35]+sumram[132][36]+sumram[132][37]+sumram[132][38]+sumram[132][39]+sumram[132][40]+sumram[132][41]+sumram[132][42]+sumram[132][43]+sumram[132][44]+sumram[132][45]+sumram[132][46]+sumram[132][47]+sumram[132][48]+sumram[132][49]+sumram[132][50]+sumram[132][51]+sumram[132][52]+sumram[132][53]+sumram[132][54]+sumram[132][55]+sumram[132][56]+sumram[132][57]+sumram[132][58]+sumram[132][59]+sumram[132][60]+sumram[132][61]+sumram[132][62]+sumram[132][63]+sumram[132][64]+sumram[132][65]+sumram[132][66]+sumram[132][67]+sumram[132][68]+sumram[132][69]+sumram[132][70]+sumram[132][71]+sumram[132][72]+sumram[132][73]+sumram[132][74]+sumram[132][75]+sumram[132][76]+sumram[132][77]+sumram[132][78]+sumram[132][79]+sumram[132][80]+sumram[132][81]+sumram[132][82]+sumram[132][83]+sumram[132][84]+sumram[132][85]+sumram[132][86]+sumram[132][87]+sumram[132][88]+sumram[132][89]+sumram[132][90]+sumram[132][91]+sumram[132][92]+sumram[132][93]+sumram[132][94]+sumram[132][95]+sumram[132][96]+sumram[132][97]+sumram[132][98]+sumram[132][99]+sumram[132][100]+sumram[132][101]+sumram[132][102]+sumram[132][103]+sumram[132][104]+sumram[132][105]+sumram[132][106]+sumram[132][107]+sumram[132][108]+sumram[132][109]+sumram[132][110]+sumram[132][111]+sumram[132][112]+sumram[132][113]+sumram[132][114]+sumram[132][115]+sumram[132][116]+sumram[132][117]+sumram[132][118]+sumram[132][119]+sumram[132][120]+sumram[132][121]+sumram[132][122]+sumram[132][123]+sumram[132][124]+sumram[132][125]+sumram[132][126]+sumram[132][127]+sumram[132][128]+sumram[132][129]+sumram[132][130]+sumram[132][131]+sumram[132][132]+sumram[132][133]+sumram[132][134]+sumram[132][135]+sumram[132][136];
    assign sumcache[133]=sumram[133][0]+sumram[133][1]+sumram[133][2]+sumram[133][3]+sumram[133][4]+sumram[133][5]+sumram[133][6]+sumram[133][7]+sumram[133][8]+sumram[133][9]+sumram[133][10]+sumram[133][11]+sumram[133][12]+sumram[133][13]+sumram[133][14]+sumram[133][15]+sumram[133][16]+sumram[133][17]+sumram[133][18]+sumram[133][19]+sumram[133][20]+sumram[133][21]+sumram[133][22]+sumram[133][23]+sumram[133][24]+sumram[133][25]+sumram[133][26]+sumram[133][27]+sumram[133][28]+sumram[133][29]+sumram[133][30]+sumram[133][31]+sumram[133][32]+sumram[133][33]+sumram[133][34]+sumram[133][35]+sumram[133][36]+sumram[133][37]+sumram[133][38]+sumram[133][39]+sumram[133][40]+sumram[133][41]+sumram[133][42]+sumram[133][43]+sumram[133][44]+sumram[133][45]+sumram[133][46]+sumram[133][47]+sumram[133][48]+sumram[133][49]+sumram[133][50]+sumram[133][51]+sumram[133][52]+sumram[133][53]+sumram[133][54]+sumram[133][55]+sumram[133][56]+sumram[133][57]+sumram[133][58]+sumram[133][59]+sumram[133][60]+sumram[133][61]+sumram[133][62]+sumram[133][63]+sumram[133][64]+sumram[133][65]+sumram[133][66]+sumram[133][67]+sumram[133][68]+sumram[133][69]+sumram[133][70]+sumram[133][71]+sumram[133][72]+sumram[133][73]+sumram[133][74]+sumram[133][75]+sumram[133][76]+sumram[133][77]+sumram[133][78]+sumram[133][79]+sumram[133][80]+sumram[133][81]+sumram[133][82]+sumram[133][83]+sumram[133][84]+sumram[133][85]+sumram[133][86]+sumram[133][87]+sumram[133][88]+sumram[133][89]+sumram[133][90]+sumram[133][91]+sumram[133][92]+sumram[133][93]+sumram[133][94]+sumram[133][95]+sumram[133][96]+sumram[133][97]+sumram[133][98]+sumram[133][99]+sumram[133][100]+sumram[133][101]+sumram[133][102]+sumram[133][103]+sumram[133][104]+sumram[133][105]+sumram[133][106]+sumram[133][107]+sumram[133][108]+sumram[133][109]+sumram[133][110]+sumram[133][111]+sumram[133][112]+sumram[133][113]+sumram[133][114]+sumram[133][115]+sumram[133][116]+sumram[133][117]+sumram[133][118]+sumram[133][119]+sumram[133][120]+sumram[133][121]+sumram[133][122]+sumram[133][123]+sumram[133][124]+sumram[133][125]+sumram[133][126]+sumram[133][127]+sumram[133][128]+sumram[133][129]+sumram[133][130]+sumram[133][131]+sumram[133][132]+sumram[133][133]+sumram[133][134]+sumram[133][135]+sumram[133][136];
    assign sumcache[134]=sumram[134][0]+sumram[134][1]+sumram[134][2]+sumram[134][3]+sumram[134][4]+sumram[134][5]+sumram[134][6]+sumram[134][7]+sumram[134][8]+sumram[134][9]+sumram[134][10]+sumram[134][11]+sumram[134][12]+sumram[134][13]+sumram[134][14]+sumram[134][15]+sumram[134][16]+sumram[134][17]+sumram[134][18]+sumram[134][19]+sumram[134][20]+sumram[134][21]+sumram[134][22]+sumram[134][23]+sumram[134][24]+sumram[134][25]+sumram[134][26]+sumram[134][27]+sumram[134][28]+sumram[134][29]+sumram[134][30]+sumram[134][31]+sumram[134][32]+sumram[134][33]+sumram[134][34]+sumram[134][35]+sumram[134][36]+sumram[134][37]+sumram[134][38]+sumram[134][39]+sumram[134][40]+sumram[134][41]+sumram[134][42]+sumram[134][43]+sumram[134][44]+sumram[134][45]+sumram[134][46]+sumram[134][47]+sumram[134][48]+sumram[134][49]+sumram[134][50]+sumram[134][51]+sumram[134][52]+sumram[134][53]+sumram[134][54]+sumram[134][55]+sumram[134][56]+sumram[134][57]+sumram[134][58]+sumram[134][59]+sumram[134][60]+sumram[134][61]+sumram[134][62]+sumram[134][63]+sumram[134][64]+sumram[134][65]+sumram[134][66]+sumram[134][67]+sumram[134][68]+sumram[134][69]+sumram[134][70]+sumram[134][71]+sumram[134][72]+sumram[134][73]+sumram[134][74]+sumram[134][75]+sumram[134][76]+sumram[134][77]+sumram[134][78]+sumram[134][79]+sumram[134][80]+sumram[134][81]+sumram[134][82]+sumram[134][83]+sumram[134][84]+sumram[134][85]+sumram[134][86]+sumram[134][87]+sumram[134][88]+sumram[134][89]+sumram[134][90]+sumram[134][91]+sumram[134][92]+sumram[134][93]+sumram[134][94]+sumram[134][95]+sumram[134][96]+sumram[134][97]+sumram[134][98]+sumram[134][99]+sumram[134][100]+sumram[134][101]+sumram[134][102]+sumram[134][103]+sumram[134][104]+sumram[134][105]+sumram[134][106]+sumram[134][107]+sumram[134][108]+sumram[134][109]+sumram[134][110]+sumram[134][111]+sumram[134][112]+sumram[134][113]+sumram[134][114]+sumram[134][115]+sumram[134][116]+sumram[134][117]+sumram[134][118]+sumram[134][119]+sumram[134][120]+sumram[134][121]+sumram[134][122]+sumram[134][123]+sumram[134][124]+sumram[134][125]+sumram[134][126]+sumram[134][127]+sumram[134][128]+sumram[134][129]+sumram[134][130]+sumram[134][131]+sumram[134][132]+sumram[134][133]+sumram[134][134]+sumram[134][135]+sumram[134][136];
    assign sumcache[135]=sumram[135][0]+sumram[135][1]+sumram[135][2]+sumram[135][3]+sumram[135][4]+sumram[135][5]+sumram[135][6]+sumram[135][7]+sumram[135][8]+sumram[135][9]+sumram[135][10]+sumram[135][11]+sumram[135][12]+sumram[135][13]+sumram[135][14]+sumram[135][15]+sumram[135][16]+sumram[135][17]+sumram[135][18]+sumram[135][19]+sumram[135][20]+sumram[135][21]+sumram[135][22]+sumram[135][23]+sumram[135][24]+sumram[135][25]+sumram[135][26]+sumram[135][27]+sumram[135][28]+sumram[135][29]+sumram[135][30]+sumram[135][31]+sumram[135][32]+sumram[135][33]+sumram[135][34]+sumram[135][35]+sumram[135][36]+sumram[135][37]+sumram[135][38]+sumram[135][39]+sumram[135][40]+sumram[135][41]+sumram[135][42]+sumram[135][43]+sumram[135][44]+sumram[135][45]+sumram[135][46]+sumram[135][47]+sumram[135][48]+sumram[135][49]+sumram[135][50]+sumram[135][51]+sumram[135][52]+sumram[135][53]+sumram[135][54]+sumram[135][55]+sumram[135][56]+sumram[135][57]+sumram[135][58]+sumram[135][59]+sumram[135][60]+sumram[135][61]+sumram[135][62]+sumram[135][63]+sumram[135][64]+sumram[135][65]+sumram[135][66]+sumram[135][67]+sumram[135][68]+sumram[135][69]+sumram[135][70]+sumram[135][71]+sumram[135][72]+sumram[135][73]+sumram[135][74]+sumram[135][75]+sumram[135][76]+sumram[135][77]+sumram[135][78]+sumram[135][79]+sumram[135][80]+sumram[135][81]+sumram[135][82]+sumram[135][83]+sumram[135][84]+sumram[135][85]+sumram[135][86]+sumram[135][87]+sumram[135][88]+sumram[135][89]+sumram[135][90]+sumram[135][91]+sumram[135][92]+sumram[135][93]+sumram[135][94]+sumram[135][95]+sumram[135][96]+sumram[135][97]+sumram[135][98]+sumram[135][99]+sumram[135][100]+sumram[135][101]+sumram[135][102]+sumram[135][103]+sumram[135][104]+sumram[135][105]+sumram[135][106]+sumram[135][107]+sumram[135][108]+sumram[135][109]+sumram[135][110]+sumram[135][111]+sumram[135][112]+sumram[135][113]+sumram[135][114]+sumram[135][115]+sumram[135][116]+sumram[135][117]+sumram[135][118]+sumram[135][119]+sumram[135][120]+sumram[135][121]+sumram[135][122]+sumram[135][123]+sumram[135][124]+sumram[135][125]+sumram[135][126]+sumram[135][127]+sumram[135][128]+sumram[135][129]+sumram[135][130]+sumram[135][131]+sumram[135][132]+sumram[135][133]+sumram[135][134]+sumram[135][135]+sumram[135][136];
    assign sumcache[136]=sumram[136][0]+sumram[136][1]+sumram[136][2]+sumram[136][3]+sumram[136][4]+sumram[136][5]+sumram[136][6]+sumram[136][7]+sumram[136][8]+sumram[136][9]+sumram[136][10]+sumram[136][11]+sumram[136][12]+sumram[136][13]+sumram[136][14]+sumram[136][15]+sumram[136][16]+sumram[136][17]+sumram[136][18]+sumram[136][19]+sumram[136][20]+sumram[136][21]+sumram[136][22]+sumram[136][23]+sumram[136][24]+sumram[136][25]+sumram[136][26]+sumram[136][27]+sumram[136][28]+sumram[136][29]+sumram[136][30]+sumram[136][31]+sumram[136][32]+sumram[136][33]+sumram[136][34]+sumram[136][35]+sumram[136][36]+sumram[136][37]+sumram[136][38]+sumram[136][39]+sumram[136][40]+sumram[136][41]+sumram[136][42]+sumram[136][43]+sumram[136][44]+sumram[136][45]+sumram[136][46]+sumram[136][47]+sumram[136][48]+sumram[136][49]+sumram[136][50]+sumram[136][51]+sumram[136][52]+sumram[136][53]+sumram[136][54]+sumram[136][55]+sumram[136][56]+sumram[136][57]+sumram[136][58]+sumram[136][59]+sumram[136][60]+sumram[136][61]+sumram[136][62]+sumram[136][63]+sumram[136][64]+sumram[136][65]+sumram[136][66]+sumram[136][67]+sumram[136][68]+sumram[136][69]+sumram[136][70]+sumram[136][71]+sumram[136][72]+sumram[136][73]+sumram[136][74]+sumram[136][75]+sumram[136][76]+sumram[136][77]+sumram[136][78]+sumram[136][79]+sumram[136][80]+sumram[136][81]+sumram[136][82]+sumram[136][83]+sumram[136][84]+sumram[136][85]+sumram[136][86]+sumram[136][87]+sumram[136][88]+sumram[136][89]+sumram[136][90]+sumram[136][91]+sumram[136][92]+sumram[136][93]+sumram[136][94]+sumram[136][95]+sumram[136][96]+sumram[136][97]+sumram[136][98]+sumram[136][99]+sumram[136][100]+sumram[136][101]+sumram[136][102]+sumram[136][103]+sumram[136][104]+sumram[136][105]+sumram[136][106]+sumram[136][107]+sumram[136][108]+sumram[136][109]+sumram[136][110]+sumram[136][111]+sumram[136][112]+sumram[136][113]+sumram[136][114]+sumram[136][115]+sumram[136][116]+sumram[136][117]+sumram[136][118]+sumram[136][119]+sumram[136][120]+sumram[136][121]+sumram[136][122]+sumram[136][123]+sumram[136][124]+sumram[136][125]+sumram[136][126]+sumram[136][127]+sumram[136][128]+sumram[136][129]+sumram[136][130]+sumram[136][131]+sumram[136][132]+sumram[136][133]+sumram[136][134]+sumram[136][135]+sumram[136][136];
    
    wire [31:0]sum_cache;
    assign sum_cache=sumcache[0]+sumcache[1]+sumcache[2]+sumcache[3]+sumcache[4]+sumcache[5]+sumcache[6]+sumcache[7]+sumcache[8]+sumcache[9]+sumcache[10]+sumcache[11]+sumcache[12]+sumcache[13]+sumcache[14]+sumcache[15]+sumcache[16]+sumcache[17]+sumcache[18]+sumcache[19]+sumcache[20]+sumcache[21]+sumcache[22]+sumcache[23]+sumcache[24]+sumcache[25]+sumcache[26]+sumcache[27]+sumcache[28]+sumcache[29]+sumcache[30]+sumcache[31]+sumcache[32]+sumcache[33]+sumcache[34]+sumcache[35]+sumcache[36]+sumcache[37]+sumcache[38]+sumcache[39]+sumcache[40]+sumcache[41]+sumcache[42]+sumcache[43]+sumcache[44]+sumcache[45]+sumcache[46]+sumcache[47]+sumcache[48]+sumcache[49]+sumcache[50]+sumcache[51]+sumcache[52]+sumcache[53]+sumcache[54]+sumcache[55]+sumcache[56]+sumcache[57]+sumcache[58]+sumcache[59]+sumcache[60]+sumcache[61]+sumcache[62]+sumcache[63]+sumcache[64]+sumcache[65]+sumcache[66]+sumcache[67]+sumcache[68]+sumcache[69]+sumcache[70]+sumcache[71]+sumcache[72]+sumcache[73]+sumcache[74]+sumcache[75]+sumcache[76]+sumcache[77]+sumcache[78]+sumcache[79]+sumcache[80]+sumcache[81]+sumcache[82]+sumcache[83]+sumcache[84]+sumcache[85]+sumcache[86]+sumcache[87]+sumcache[88]+sumcache[89]+sumcache[90]+sumcache[91]+sumcache[92]+sumcache[93]+sumcache[94]+sumcache[95]+sumcache[96]+sumcache[97]+sumcache[98]+sumcache[99]+sumcache[100]+sumcache[101]+sumcache[102]+sumcache[103]+sumcache[104]+sumcache[105]+sumcache[106]+sumcache[107]+sumcache[108]+sumcache[109]+sumcache[110]+sumcache[111]+sumcache[112]+sumcache[113]+sumcache[114]+sumcache[115]+sumcache[116]+sumcache[117]+sumcache[118]+sumcache[119]+sumcache[120]+sumcache[121]+sumcache[122]+sumcache[123]+sumcache[124]+sumcache[125]+sumcache[126]+sumcache[127]+sumcache[128]+sumcache[129]+sumcache[130]+sumcache[131]+sumcache[132]+sumcache[133]+sumcache[134]+sumcache[135]+sumcache[136];
    
    genvar a,b;
    generate
        for (a=0;a<size;a=a+1)
        begin: ram_row
            for (b=0;b<size;b=b+1)
            begin: ram_column
                always @(posedge clk) ram[a][b]<=ram[a][b]-sumram[a][b];
            end    
        end
    endgenerate
    
    always @(posedge clk)
    begin
        if(rst)sum<=0;
        else sum<=sum+sum_cache;
    end
    
endmodule

