`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.01.2026 18:58:52
// Design Name: 
// Module Name: Main
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Main(
    input clk,rst,
    output reg [63:0]ans1,ans2
    );
    parameter size=141;
    
    reg [size-1:0]ram[size/2-1:0];
    reg [63:0]ans2_ram[size-1:0];
    initial 
    begin
        ram[0][0]=0;ram[0][1]=0;ram[0][2]=0;ram[0][3]=0;ram[0][4]=0;ram[0][5]=0;ram[0][6]=0;ram[0][7]=0;ram[0][8]=0;ram[0][9]=0;ram[0][10]=0;ram[0][11]=0;ram[0][12]=0;ram[0][13]=0;ram[0][14]=0;ram[0][15]=0;ram[0][16]=0;ram[0][17]=0;ram[0][18]=0;ram[0][19]=0;ram[0][20]=0;ram[0][21]=0;ram[0][22]=0;ram[0][23]=0;ram[0][24]=0;ram[0][25]=0;ram[0][26]=0;ram[0][27]=0;ram[0][28]=0;ram[0][29]=0;ram[0][30]=0;ram[0][31]=0;ram[0][32]=0;ram[0][33]=0;ram[0][34]=0;ram[0][35]=0;ram[0][36]=0;ram[0][37]=0;ram[0][38]=0;ram[0][39]=0;ram[0][40]=0;ram[0][41]=0;ram[0][42]=0;ram[0][43]=0;ram[0][44]=0;ram[0][45]=0;ram[0][46]=0;ram[0][47]=0;ram[0][48]=0;ram[0][49]=0;ram[0][50]=0;ram[0][51]=0;ram[0][52]=0;ram[0][53]=0;ram[0][54]=0;ram[0][55]=0;ram[0][56]=0;ram[0][57]=0;ram[0][58]=0;ram[0][59]=0;ram[0][60]=0;ram[0][61]=0;ram[0][62]=0;ram[0][63]=0;ram[0][64]=0;ram[0][65]=0;ram[0][66]=0;ram[0][67]=0;ram[0][68]=0;ram[0][69]=0;ram[0][70]=1;ram[0][71]=0;ram[0][72]=0;ram[0][73]=0;ram[0][74]=0;ram[0][75]=0;ram[0][76]=0;ram[0][77]=0;ram[0][78]=0;ram[0][79]=0;ram[0][80]=0;ram[0][81]=0;ram[0][82]=0;ram[0][83]=0;ram[0][84]=0;ram[0][85]=0;ram[0][86]=0;ram[0][87]=0;ram[0][88]=0;ram[0][89]=0;ram[0][90]=0;ram[0][91]=0;ram[0][92]=0;ram[0][93]=0;ram[0][94]=0;ram[0][95]=0;ram[0][96]=0;ram[0][97]=0;ram[0][98]=0;ram[0][99]=0;ram[0][100]=0;ram[0][101]=0;ram[0][102]=0;ram[0][103]=0;ram[0][104]=0;ram[0][105]=0;ram[0][106]=0;ram[0][107]=0;ram[0][108]=0;ram[0][109]=0;ram[0][110]=0;ram[0][111]=0;ram[0][112]=0;ram[0][113]=0;ram[0][114]=0;ram[0][115]=0;ram[0][116]=0;ram[0][117]=0;ram[0][118]=0;ram[0][119]=0;ram[0][120]=0;ram[0][121]=0;ram[0][122]=0;ram[0][123]=0;ram[0][124]=0;ram[0][125]=0;ram[0][126]=0;ram[0][127]=0;ram[0][128]=0;ram[0][129]=0;ram[0][130]=0;ram[0][131]=0;ram[0][132]=0;ram[0][133]=0;ram[0][134]=0;ram[0][135]=0;ram[0][136]=0;ram[0][137]=0;ram[0][138]=0;ram[0][139]=0;ram[0][140]=0;
        ram[1][0]=0;ram[1][1]=0;ram[1][2]=0;ram[1][3]=0;ram[1][4]=0;ram[1][5]=0;ram[1][6]=0;ram[1][7]=0;ram[1][8]=0;ram[1][9]=0;ram[1][10]=0;ram[1][11]=0;ram[1][12]=0;ram[1][13]=0;ram[1][14]=0;ram[1][15]=0;ram[1][16]=0;ram[1][17]=0;ram[1][18]=0;ram[1][19]=0;ram[1][20]=0;ram[1][21]=0;ram[1][22]=0;ram[1][23]=0;ram[1][24]=0;ram[1][25]=0;ram[1][26]=0;ram[1][27]=0;ram[1][28]=0;ram[1][29]=0;ram[1][30]=0;ram[1][31]=0;ram[1][32]=0;ram[1][33]=0;ram[1][34]=0;ram[1][35]=0;ram[1][36]=0;ram[1][37]=0;ram[1][38]=0;ram[1][39]=0;ram[1][40]=0;ram[1][41]=0;ram[1][42]=0;ram[1][43]=0;ram[1][44]=0;ram[1][45]=0;ram[1][46]=0;ram[1][47]=0;ram[1][48]=0;ram[1][49]=0;ram[1][50]=0;ram[1][51]=0;ram[1][52]=0;ram[1][53]=0;ram[1][54]=0;ram[1][55]=0;ram[1][56]=0;ram[1][57]=0;ram[1][58]=0;ram[1][59]=0;ram[1][60]=0;ram[1][61]=0;ram[1][62]=0;ram[1][63]=0;ram[1][64]=0;ram[1][65]=0;ram[1][66]=0;ram[1][67]=0;ram[1][68]=0;ram[1][69]=1;ram[1][70]=0;ram[1][71]=1;ram[1][72]=0;ram[1][73]=0;ram[1][74]=0;ram[1][75]=0;ram[1][76]=0;ram[1][77]=0;ram[1][78]=0;ram[1][79]=0;ram[1][80]=0;ram[1][81]=0;ram[1][82]=0;ram[1][83]=0;ram[1][84]=0;ram[1][85]=0;ram[1][86]=0;ram[1][87]=0;ram[1][88]=0;ram[1][89]=0;ram[1][90]=0;ram[1][91]=0;ram[1][92]=0;ram[1][93]=0;ram[1][94]=0;ram[1][95]=0;ram[1][96]=0;ram[1][97]=0;ram[1][98]=0;ram[1][99]=0;ram[1][100]=0;ram[1][101]=0;ram[1][102]=0;ram[1][103]=0;ram[1][104]=0;ram[1][105]=0;ram[1][106]=0;ram[1][107]=0;ram[1][108]=0;ram[1][109]=0;ram[1][110]=0;ram[1][111]=0;ram[1][112]=0;ram[1][113]=0;ram[1][114]=0;ram[1][115]=0;ram[1][116]=0;ram[1][117]=0;ram[1][118]=0;ram[1][119]=0;ram[1][120]=0;ram[1][121]=0;ram[1][122]=0;ram[1][123]=0;ram[1][124]=0;ram[1][125]=0;ram[1][126]=0;ram[1][127]=0;ram[1][128]=0;ram[1][129]=0;ram[1][130]=0;ram[1][131]=0;ram[1][132]=0;ram[1][133]=0;ram[1][134]=0;ram[1][135]=0;ram[1][136]=0;ram[1][137]=0;ram[1][138]=0;ram[1][139]=0;ram[1][140]=0;
        ram[2][0]=0;ram[2][1]=0;ram[2][2]=0;ram[2][3]=0;ram[2][4]=0;ram[2][5]=0;ram[2][6]=0;ram[2][7]=0;ram[2][8]=0;ram[2][9]=0;ram[2][10]=0;ram[2][11]=0;ram[2][12]=0;ram[2][13]=0;ram[2][14]=0;ram[2][15]=0;ram[2][16]=0;ram[2][17]=0;ram[2][18]=0;ram[2][19]=0;ram[2][20]=0;ram[2][21]=0;ram[2][22]=0;ram[2][23]=0;ram[2][24]=0;ram[2][25]=0;ram[2][26]=0;ram[2][27]=0;ram[2][28]=0;ram[2][29]=0;ram[2][30]=0;ram[2][31]=0;ram[2][32]=0;ram[2][33]=0;ram[2][34]=0;ram[2][35]=0;ram[2][36]=0;ram[2][37]=0;ram[2][38]=0;ram[2][39]=0;ram[2][40]=0;ram[2][41]=0;ram[2][42]=0;ram[2][43]=0;ram[2][44]=0;ram[2][45]=0;ram[2][46]=0;ram[2][47]=0;ram[2][48]=0;ram[2][49]=0;ram[2][50]=0;ram[2][51]=0;ram[2][52]=0;ram[2][53]=0;ram[2][54]=0;ram[2][55]=0;ram[2][56]=0;ram[2][57]=0;ram[2][58]=0;ram[2][59]=0;ram[2][60]=0;ram[2][61]=0;ram[2][62]=0;ram[2][63]=0;ram[2][64]=0;ram[2][65]=0;ram[2][66]=0;ram[2][67]=0;ram[2][68]=1;ram[2][69]=0;ram[2][70]=0;ram[2][71]=0;ram[2][72]=1;ram[2][73]=0;ram[2][74]=0;ram[2][75]=0;ram[2][76]=0;ram[2][77]=0;ram[2][78]=0;ram[2][79]=0;ram[2][80]=0;ram[2][81]=0;ram[2][82]=0;ram[2][83]=0;ram[2][84]=0;ram[2][85]=0;ram[2][86]=0;ram[2][87]=0;ram[2][88]=0;ram[2][89]=0;ram[2][90]=0;ram[2][91]=0;ram[2][92]=0;ram[2][93]=0;ram[2][94]=0;ram[2][95]=0;ram[2][96]=0;ram[2][97]=0;ram[2][98]=0;ram[2][99]=0;ram[2][100]=0;ram[2][101]=0;ram[2][102]=0;ram[2][103]=0;ram[2][104]=0;ram[2][105]=0;ram[2][106]=0;ram[2][107]=0;ram[2][108]=0;ram[2][109]=0;ram[2][110]=0;ram[2][111]=0;ram[2][112]=0;ram[2][113]=0;ram[2][114]=0;ram[2][115]=0;ram[2][116]=0;ram[2][117]=0;ram[2][118]=0;ram[2][119]=0;ram[2][120]=0;ram[2][121]=0;ram[2][122]=0;ram[2][123]=0;ram[2][124]=0;ram[2][125]=0;ram[2][126]=0;ram[2][127]=0;ram[2][128]=0;ram[2][129]=0;ram[2][130]=0;ram[2][131]=0;ram[2][132]=0;ram[2][133]=0;ram[2][134]=0;ram[2][135]=0;ram[2][136]=0;ram[2][137]=0;ram[2][138]=0;ram[2][139]=0;ram[2][140]=0;
        ram[3][0]=0;ram[3][1]=0;ram[3][2]=0;ram[3][3]=0;ram[3][4]=0;ram[3][5]=0;ram[3][6]=0;ram[3][7]=0;ram[3][8]=0;ram[3][9]=0;ram[3][10]=0;ram[3][11]=0;ram[3][12]=0;ram[3][13]=0;ram[3][14]=0;ram[3][15]=0;ram[3][16]=0;ram[3][17]=0;ram[3][18]=0;ram[3][19]=0;ram[3][20]=0;ram[3][21]=0;ram[3][22]=0;ram[3][23]=0;ram[3][24]=0;ram[3][25]=0;ram[3][26]=0;ram[3][27]=0;ram[3][28]=0;ram[3][29]=0;ram[3][30]=0;ram[3][31]=0;ram[3][32]=0;ram[3][33]=0;ram[3][34]=0;ram[3][35]=0;ram[3][36]=0;ram[3][37]=0;ram[3][38]=0;ram[3][39]=0;ram[3][40]=0;ram[3][41]=0;ram[3][42]=0;ram[3][43]=0;ram[3][44]=0;ram[3][45]=0;ram[3][46]=0;ram[3][47]=0;ram[3][48]=0;ram[3][49]=0;ram[3][50]=0;ram[3][51]=0;ram[3][52]=0;ram[3][53]=0;ram[3][54]=0;ram[3][55]=0;ram[3][56]=0;ram[3][57]=0;ram[3][58]=0;ram[3][59]=0;ram[3][60]=0;ram[3][61]=0;ram[3][62]=0;ram[3][63]=0;ram[3][64]=0;ram[3][65]=0;ram[3][66]=0;ram[3][67]=1;ram[3][68]=0;ram[3][69]=0;ram[3][70]=0;ram[3][71]=1;ram[3][72]=0;ram[3][73]=1;ram[3][74]=0;ram[3][75]=0;ram[3][76]=0;ram[3][77]=0;ram[3][78]=0;ram[3][79]=0;ram[3][80]=0;ram[3][81]=0;ram[3][82]=0;ram[3][83]=0;ram[3][84]=0;ram[3][85]=0;ram[3][86]=0;ram[3][87]=0;ram[3][88]=0;ram[3][89]=0;ram[3][90]=0;ram[3][91]=0;ram[3][92]=0;ram[3][93]=0;ram[3][94]=0;ram[3][95]=0;ram[3][96]=0;ram[3][97]=0;ram[3][98]=0;ram[3][99]=0;ram[3][100]=0;ram[3][101]=0;ram[3][102]=0;ram[3][103]=0;ram[3][104]=0;ram[3][105]=0;ram[3][106]=0;ram[3][107]=0;ram[3][108]=0;ram[3][109]=0;ram[3][110]=0;ram[3][111]=0;ram[3][112]=0;ram[3][113]=0;ram[3][114]=0;ram[3][115]=0;ram[3][116]=0;ram[3][117]=0;ram[3][118]=0;ram[3][119]=0;ram[3][120]=0;ram[3][121]=0;ram[3][122]=0;ram[3][123]=0;ram[3][124]=0;ram[3][125]=0;ram[3][126]=0;ram[3][127]=0;ram[3][128]=0;ram[3][129]=0;ram[3][130]=0;ram[3][131]=0;ram[3][132]=0;ram[3][133]=0;ram[3][134]=0;ram[3][135]=0;ram[3][136]=0;ram[3][137]=0;ram[3][138]=0;ram[3][139]=0;ram[3][140]=0;
        ram[4][0]=0;ram[4][1]=0;ram[4][2]=0;ram[4][3]=0;ram[4][4]=0;ram[4][5]=0;ram[4][6]=0;ram[4][7]=0;ram[4][8]=0;ram[4][9]=0;ram[4][10]=0;ram[4][11]=0;ram[4][12]=0;ram[4][13]=0;ram[4][14]=0;ram[4][15]=0;ram[4][16]=0;ram[4][17]=0;ram[4][18]=0;ram[4][19]=0;ram[4][20]=0;ram[4][21]=0;ram[4][22]=0;ram[4][23]=0;ram[4][24]=0;ram[4][25]=0;ram[4][26]=0;ram[4][27]=0;ram[4][28]=0;ram[4][29]=0;ram[4][30]=0;ram[4][31]=0;ram[4][32]=0;ram[4][33]=0;ram[4][34]=0;ram[4][35]=0;ram[4][36]=0;ram[4][37]=0;ram[4][38]=0;ram[4][39]=0;ram[4][40]=0;ram[4][41]=0;ram[4][42]=0;ram[4][43]=0;ram[4][44]=0;ram[4][45]=0;ram[4][46]=0;ram[4][47]=0;ram[4][48]=0;ram[4][49]=0;ram[4][50]=0;ram[4][51]=0;ram[4][52]=0;ram[4][53]=0;ram[4][54]=0;ram[4][55]=0;ram[4][56]=0;ram[4][57]=0;ram[4][58]=0;ram[4][59]=0;ram[4][60]=0;ram[4][61]=0;ram[4][62]=0;ram[4][63]=0;ram[4][64]=0;ram[4][65]=0;ram[4][66]=1;ram[4][67]=0;ram[4][68]=1;ram[4][69]=0;ram[4][70]=0;ram[4][71]=0;ram[4][72]=1;ram[4][73]=0;ram[4][74]=1;ram[4][75]=0;ram[4][76]=0;ram[4][77]=0;ram[4][78]=0;ram[4][79]=0;ram[4][80]=0;ram[4][81]=0;ram[4][82]=0;ram[4][83]=0;ram[4][84]=0;ram[4][85]=0;ram[4][86]=0;ram[4][87]=0;ram[4][88]=0;ram[4][89]=0;ram[4][90]=0;ram[4][91]=0;ram[4][92]=0;ram[4][93]=0;ram[4][94]=0;ram[4][95]=0;ram[4][96]=0;ram[4][97]=0;ram[4][98]=0;ram[4][99]=0;ram[4][100]=0;ram[4][101]=0;ram[4][102]=0;ram[4][103]=0;ram[4][104]=0;ram[4][105]=0;ram[4][106]=0;ram[4][107]=0;ram[4][108]=0;ram[4][109]=0;ram[4][110]=0;ram[4][111]=0;ram[4][112]=0;ram[4][113]=0;ram[4][114]=0;ram[4][115]=0;ram[4][116]=0;ram[4][117]=0;ram[4][118]=0;ram[4][119]=0;ram[4][120]=0;ram[4][121]=0;ram[4][122]=0;ram[4][123]=0;ram[4][124]=0;ram[4][125]=0;ram[4][126]=0;ram[4][127]=0;ram[4][128]=0;ram[4][129]=0;ram[4][130]=0;ram[4][131]=0;ram[4][132]=0;ram[4][133]=0;ram[4][134]=0;ram[4][135]=0;ram[4][136]=0;ram[4][137]=0;ram[4][138]=0;ram[4][139]=0;ram[4][140]=0;
        ram[5][0]=0;ram[5][1]=0;ram[5][2]=0;ram[5][3]=0;ram[5][4]=0;ram[5][5]=0;ram[5][6]=0;ram[5][7]=0;ram[5][8]=0;ram[5][9]=0;ram[5][10]=0;ram[5][11]=0;ram[5][12]=0;ram[5][13]=0;ram[5][14]=0;ram[5][15]=0;ram[5][16]=0;ram[5][17]=0;ram[5][18]=0;ram[5][19]=0;ram[5][20]=0;ram[5][21]=0;ram[5][22]=0;ram[5][23]=0;ram[5][24]=0;ram[5][25]=0;ram[5][26]=0;ram[5][27]=0;ram[5][28]=0;ram[5][29]=0;ram[5][30]=0;ram[5][31]=0;ram[5][32]=0;ram[5][33]=0;ram[5][34]=0;ram[5][35]=0;ram[5][36]=0;ram[5][37]=0;ram[5][38]=0;ram[5][39]=0;ram[5][40]=0;ram[5][41]=0;ram[5][42]=0;ram[5][43]=0;ram[5][44]=0;ram[5][45]=0;ram[5][46]=0;ram[5][47]=0;ram[5][48]=0;ram[5][49]=0;ram[5][50]=0;ram[5][51]=0;ram[5][52]=0;ram[5][53]=0;ram[5][54]=0;ram[5][55]=0;ram[5][56]=0;ram[5][57]=0;ram[5][58]=0;ram[5][59]=0;ram[5][60]=0;ram[5][61]=0;ram[5][62]=0;ram[5][63]=0;ram[5][64]=0;ram[5][65]=1;ram[5][66]=0;ram[5][67]=1;ram[5][68]=0;ram[5][69]=1;ram[5][70]=0;ram[5][71]=1;ram[5][72]=0;ram[5][73]=1;ram[5][74]=0;ram[5][75]=1;ram[5][76]=0;ram[5][77]=0;ram[5][78]=0;ram[5][79]=0;ram[5][80]=0;ram[5][81]=0;ram[5][82]=0;ram[5][83]=0;ram[5][84]=0;ram[5][85]=0;ram[5][86]=0;ram[5][87]=0;ram[5][88]=0;ram[5][89]=0;ram[5][90]=0;ram[5][91]=0;ram[5][92]=0;ram[5][93]=0;ram[5][94]=0;ram[5][95]=0;ram[5][96]=0;ram[5][97]=0;ram[5][98]=0;ram[5][99]=0;ram[5][100]=0;ram[5][101]=0;ram[5][102]=0;ram[5][103]=0;ram[5][104]=0;ram[5][105]=0;ram[5][106]=0;ram[5][107]=0;ram[5][108]=0;ram[5][109]=0;ram[5][110]=0;ram[5][111]=0;ram[5][112]=0;ram[5][113]=0;ram[5][114]=0;ram[5][115]=0;ram[5][116]=0;ram[5][117]=0;ram[5][118]=0;ram[5][119]=0;ram[5][120]=0;ram[5][121]=0;ram[5][122]=0;ram[5][123]=0;ram[5][124]=0;ram[5][125]=0;ram[5][126]=0;ram[5][127]=0;ram[5][128]=0;ram[5][129]=0;ram[5][130]=0;ram[5][131]=0;ram[5][132]=0;ram[5][133]=0;ram[5][134]=0;ram[5][135]=0;ram[5][136]=0;ram[5][137]=0;ram[5][138]=0;ram[5][139]=0;ram[5][140]=0;
        ram[6][0]=0;ram[6][1]=0;ram[6][2]=0;ram[6][3]=0;ram[6][4]=0;ram[6][5]=0;ram[6][6]=0;ram[6][7]=0;ram[6][8]=0;ram[6][9]=0;ram[6][10]=0;ram[6][11]=0;ram[6][12]=0;ram[6][13]=0;ram[6][14]=0;ram[6][15]=0;ram[6][16]=0;ram[6][17]=0;ram[6][18]=0;ram[6][19]=0;ram[6][20]=0;ram[6][21]=0;ram[6][22]=0;ram[6][23]=0;ram[6][24]=0;ram[6][25]=0;ram[6][26]=0;ram[6][27]=0;ram[6][28]=0;ram[6][29]=0;ram[6][30]=0;ram[6][31]=0;ram[6][32]=0;ram[6][33]=0;ram[6][34]=0;ram[6][35]=0;ram[6][36]=0;ram[6][37]=0;ram[6][38]=0;ram[6][39]=0;ram[6][40]=0;ram[6][41]=0;ram[6][42]=0;ram[6][43]=0;ram[6][44]=0;ram[6][45]=0;ram[6][46]=0;ram[6][47]=0;ram[6][48]=0;ram[6][49]=0;ram[6][50]=0;ram[6][51]=0;ram[6][52]=0;ram[6][53]=0;ram[6][54]=0;ram[6][55]=0;ram[6][56]=0;ram[6][57]=0;ram[6][58]=0;ram[6][59]=0;ram[6][60]=0;ram[6][61]=0;ram[6][62]=0;ram[6][63]=0;ram[6][64]=1;ram[6][65]=0;ram[6][66]=1;ram[6][67]=0;ram[6][68]=0;ram[6][69]=0;ram[6][70]=1;ram[6][71]=0;ram[6][72]=0;ram[6][73]=0;ram[6][74]=1;ram[6][75]=0;ram[6][76]=1;ram[6][77]=0;ram[6][78]=0;ram[6][79]=0;ram[6][80]=0;ram[6][81]=0;ram[6][82]=0;ram[6][83]=0;ram[6][84]=0;ram[6][85]=0;ram[6][86]=0;ram[6][87]=0;ram[6][88]=0;ram[6][89]=0;ram[6][90]=0;ram[6][91]=0;ram[6][92]=0;ram[6][93]=0;ram[6][94]=0;ram[6][95]=0;ram[6][96]=0;ram[6][97]=0;ram[6][98]=0;ram[6][99]=0;ram[6][100]=0;ram[6][101]=0;ram[6][102]=0;ram[6][103]=0;ram[6][104]=0;ram[6][105]=0;ram[6][106]=0;ram[6][107]=0;ram[6][108]=0;ram[6][109]=0;ram[6][110]=0;ram[6][111]=0;ram[6][112]=0;ram[6][113]=0;ram[6][114]=0;ram[6][115]=0;ram[6][116]=0;ram[6][117]=0;ram[6][118]=0;ram[6][119]=0;ram[6][120]=0;ram[6][121]=0;ram[6][122]=0;ram[6][123]=0;ram[6][124]=0;ram[6][125]=0;ram[6][126]=0;ram[6][127]=0;ram[6][128]=0;ram[6][129]=0;ram[6][130]=0;ram[6][131]=0;ram[6][132]=0;ram[6][133]=0;ram[6][134]=0;ram[6][135]=0;ram[6][136]=0;ram[6][137]=0;ram[6][138]=0;ram[6][139]=0;ram[6][140]=0;
        ram[7][0]=0;ram[7][1]=0;ram[7][2]=0;ram[7][3]=0;ram[7][4]=0;ram[7][5]=0;ram[7][6]=0;ram[7][7]=0;ram[7][8]=0;ram[7][9]=0;ram[7][10]=0;ram[7][11]=0;ram[7][12]=0;ram[7][13]=0;ram[7][14]=0;ram[7][15]=0;ram[7][16]=0;ram[7][17]=0;ram[7][18]=0;ram[7][19]=0;ram[7][20]=0;ram[7][21]=0;ram[7][22]=0;ram[7][23]=0;ram[7][24]=0;ram[7][25]=0;ram[7][26]=0;ram[7][27]=0;ram[7][28]=0;ram[7][29]=0;ram[7][30]=0;ram[7][31]=0;ram[7][32]=0;ram[7][33]=0;ram[7][34]=0;ram[7][35]=0;ram[7][36]=0;ram[7][37]=0;ram[7][38]=0;ram[7][39]=0;ram[7][40]=0;ram[7][41]=0;ram[7][42]=0;ram[7][43]=0;ram[7][44]=0;ram[7][45]=0;ram[7][46]=0;ram[7][47]=0;ram[7][48]=0;ram[7][49]=0;ram[7][50]=0;ram[7][51]=0;ram[7][52]=0;ram[7][53]=0;ram[7][54]=0;ram[7][55]=0;ram[7][56]=0;ram[7][57]=0;ram[7][58]=0;ram[7][59]=0;ram[7][60]=0;ram[7][61]=0;ram[7][62]=0;ram[7][63]=1;ram[7][64]=0;ram[7][65]=1;ram[7][66]=0;ram[7][67]=1;ram[7][68]=0;ram[7][69]=0;ram[7][70]=0;ram[7][71]=1;ram[7][72]=0;ram[7][73]=1;ram[7][74]=0;ram[7][75]=1;ram[7][76]=0;ram[7][77]=1;ram[7][78]=0;ram[7][79]=0;ram[7][80]=0;ram[7][81]=0;ram[7][82]=0;ram[7][83]=0;ram[7][84]=0;ram[7][85]=0;ram[7][86]=0;ram[7][87]=0;ram[7][88]=0;ram[7][89]=0;ram[7][90]=0;ram[7][91]=0;ram[7][92]=0;ram[7][93]=0;ram[7][94]=0;ram[7][95]=0;ram[7][96]=0;ram[7][97]=0;ram[7][98]=0;ram[7][99]=0;ram[7][100]=0;ram[7][101]=0;ram[7][102]=0;ram[7][103]=0;ram[7][104]=0;ram[7][105]=0;ram[7][106]=0;ram[7][107]=0;ram[7][108]=0;ram[7][109]=0;ram[7][110]=0;ram[7][111]=0;ram[7][112]=0;ram[7][113]=0;ram[7][114]=0;ram[7][115]=0;ram[7][116]=0;ram[7][117]=0;ram[7][118]=0;ram[7][119]=0;ram[7][120]=0;ram[7][121]=0;ram[7][122]=0;ram[7][123]=0;ram[7][124]=0;ram[7][125]=0;ram[7][126]=0;ram[7][127]=0;ram[7][128]=0;ram[7][129]=0;ram[7][130]=0;ram[7][131]=0;ram[7][132]=0;ram[7][133]=0;ram[7][134]=0;ram[7][135]=0;ram[7][136]=0;ram[7][137]=0;ram[7][138]=0;ram[7][139]=0;ram[7][140]=0;
        ram[8][0]=0;ram[8][1]=0;ram[8][2]=0;ram[8][3]=0;ram[8][4]=0;ram[8][5]=0;ram[8][6]=0;ram[8][7]=0;ram[8][8]=0;ram[8][9]=0;ram[8][10]=0;ram[8][11]=0;ram[8][12]=0;ram[8][13]=0;ram[8][14]=0;ram[8][15]=0;ram[8][16]=0;ram[8][17]=0;ram[8][18]=0;ram[8][19]=0;ram[8][20]=0;ram[8][21]=0;ram[8][22]=0;ram[8][23]=0;ram[8][24]=0;ram[8][25]=0;ram[8][26]=0;ram[8][27]=0;ram[8][28]=0;ram[8][29]=0;ram[8][30]=0;ram[8][31]=0;ram[8][32]=0;ram[8][33]=0;ram[8][34]=0;ram[8][35]=0;ram[8][36]=0;ram[8][37]=0;ram[8][38]=0;ram[8][39]=0;ram[8][40]=0;ram[8][41]=0;ram[8][42]=0;ram[8][43]=0;ram[8][44]=0;ram[8][45]=0;ram[8][46]=0;ram[8][47]=0;ram[8][48]=0;ram[8][49]=0;ram[8][50]=0;ram[8][51]=0;ram[8][52]=0;ram[8][53]=0;ram[8][54]=0;ram[8][55]=0;ram[8][56]=0;ram[8][57]=0;ram[8][58]=0;ram[8][59]=0;ram[8][60]=0;ram[8][61]=0;ram[8][62]=1;ram[8][63]=0;ram[8][64]=0;ram[8][65]=0;ram[8][66]=1;ram[8][67]=0;ram[8][68]=1;ram[8][69]=0;ram[8][70]=0;ram[8][71]=0;ram[8][72]=0;ram[8][73]=0;ram[8][74]=1;ram[8][75]=0;ram[8][76]=1;ram[8][77]=0;ram[8][78]=1;ram[8][79]=0;ram[8][80]=0;ram[8][81]=0;ram[8][82]=0;ram[8][83]=0;ram[8][84]=0;ram[8][85]=0;ram[8][86]=0;ram[8][87]=0;ram[8][88]=0;ram[8][89]=0;ram[8][90]=0;ram[8][91]=0;ram[8][92]=0;ram[8][93]=0;ram[8][94]=0;ram[8][95]=0;ram[8][96]=0;ram[8][97]=0;ram[8][98]=0;ram[8][99]=0;ram[8][100]=0;ram[8][101]=0;ram[8][102]=0;ram[8][103]=0;ram[8][104]=0;ram[8][105]=0;ram[8][106]=0;ram[8][107]=0;ram[8][108]=0;ram[8][109]=0;ram[8][110]=0;ram[8][111]=0;ram[8][112]=0;ram[8][113]=0;ram[8][114]=0;ram[8][115]=0;ram[8][116]=0;ram[8][117]=0;ram[8][118]=0;ram[8][119]=0;ram[8][120]=0;ram[8][121]=0;ram[8][122]=0;ram[8][123]=0;ram[8][124]=0;ram[8][125]=0;ram[8][126]=0;ram[8][127]=0;ram[8][128]=0;ram[8][129]=0;ram[8][130]=0;ram[8][131]=0;ram[8][132]=0;ram[8][133]=0;ram[8][134]=0;ram[8][135]=0;ram[8][136]=0;ram[8][137]=0;ram[8][138]=0;ram[8][139]=0;ram[8][140]=0;
        ram[9][0]=0;ram[9][1]=0;ram[9][2]=0;ram[9][3]=0;ram[9][4]=0;ram[9][5]=0;ram[9][6]=0;ram[9][7]=0;ram[9][8]=0;ram[9][9]=0;ram[9][10]=0;ram[9][11]=0;ram[9][12]=0;ram[9][13]=0;ram[9][14]=0;ram[9][15]=0;ram[9][16]=0;ram[9][17]=0;ram[9][18]=0;ram[9][19]=0;ram[9][20]=0;ram[9][21]=0;ram[9][22]=0;ram[9][23]=0;ram[9][24]=0;ram[9][25]=0;ram[9][26]=0;ram[9][27]=0;ram[9][28]=0;ram[9][29]=0;ram[9][30]=0;ram[9][31]=0;ram[9][32]=0;ram[9][33]=0;ram[9][34]=0;ram[9][35]=0;ram[9][36]=0;ram[9][37]=0;ram[9][38]=0;ram[9][39]=0;ram[9][40]=0;ram[9][41]=0;ram[9][42]=0;ram[9][43]=0;ram[9][44]=0;ram[9][45]=0;ram[9][46]=0;ram[9][47]=0;ram[9][48]=0;ram[9][49]=0;ram[9][50]=0;ram[9][51]=0;ram[9][52]=0;ram[9][53]=0;ram[9][54]=0;ram[9][55]=0;ram[9][56]=0;ram[9][57]=0;ram[9][58]=0;ram[9][59]=0;ram[9][60]=0;ram[9][61]=1;ram[9][62]=0;ram[9][63]=0;ram[9][64]=0;ram[9][65]=1;ram[9][66]=0;ram[9][67]=1;ram[9][68]=0;ram[9][69]=0;ram[9][70]=0;ram[9][71]=1;ram[9][72]=0;ram[9][73]=0;ram[9][74]=0;ram[9][75]=0;ram[9][76]=0;ram[9][77]=1;ram[9][78]=0;ram[9][79]=1;ram[9][80]=0;ram[9][81]=0;ram[9][82]=0;ram[9][83]=0;ram[9][84]=0;ram[9][85]=0;ram[9][86]=0;ram[9][87]=0;ram[9][88]=0;ram[9][89]=0;ram[9][90]=0;ram[9][91]=0;ram[9][92]=0;ram[9][93]=0;ram[9][94]=0;ram[9][95]=0;ram[9][96]=0;ram[9][97]=0;ram[9][98]=0;ram[9][99]=0;ram[9][100]=0;ram[9][101]=0;ram[9][102]=0;ram[9][103]=0;ram[9][104]=0;ram[9][105]=0;ram[9][106]=0;ram[9][107]=0;ram[9][108]=0;ram[9][109]=0;ram[9][110]=0;ram[9][111]=0;ram[9][112]=0;ram[9][113]=0;ram[9][114]=0;ram[9][115]=0;ram[9][116]=0;ram[9][117]=0;ram[9][118]=0;ram[9][119]=0;ram[9][120]=0;ram[9][121]=0;ram[9][122]=0;ram[9][123]=0;ram[9][124]=0;ram[9][125]=0;ram[9][126]=0;ram[9][127]=0;ram[9][128]=0;ram[9][129]=0;ram[9][130]=0;ram[9][131]=0;ram[9][132]=0;ram[9][133]=0;ram[9][134]=0;ram[9][135]=0;ram[9][136]=0;ram[9][137]=0;ram[9][138]=0;ram[9][139]=0;ram[9][140]=0;
        ram[10][0]=0;ram[10][1]=0;ram[10][2]=0;ram[10][3]=0;ram[10][4]=0;ram[10][5]=0;ram[10][6]=0;ram[10][7]=0;ram[10][8]=0;ram[10][9]=0;ram[10][10]=0;ram[10][11]=0;ram[10][12]=0;ram[10][13]=0;ram[10][14]=0;ram[10][15]=0;ram[10][16]=0;ram[10][17]=0;ram[10][18]=0;ram[10][19]=0;ram[10][20]=0;ram[10][21]=0;ram[10][22]=0;ram[10][23]=0;ram[10][24]=0;ram[10][25]=0;ram[10][26]=0;ram[10][27]=0;ram[10][28]=0;ram[10][29]=0;ram[10][30]=0;ram[10][31]=0;ram[10][32]=0;ram[10][33]=0;ram[10][34]=0;ram[10][35]=0;ram[10][36]=0;ram[10][37]=0;ram[10][38]=0;ram[10][39]=0;ram[10][40]=0;ram[10][41]=0;ram[10][42]=0;ram[10][43]=0;ram[10][44]=0;ram[10][45]=0;ram[10][46]=0;ram[10][47]=0;ram[10][48]=0;ram[10][49]=0;ram[10][50]=0;ram[10][51]=0;ram[10][52]=0;ram[10][53]=0;ram[10][54]=0;ram[10][55]=0;ram[10][56]=0;ram[10][57]=0;ram[10][58]=0;ram[10][59]=0;ram[10][60]=1;ram[10][61]=0;ram[10][62]=1;ram[10][63]=0;ram[10][64]=0;ram[10][65]=0;ram[10][66]=0;ram[10][67]=0;ram[10][68]=1;ram[10][69]=0;ram[10][70]=1;ram[10][71]=0;ram[10][72]=1;ram[10][73]=0;ram[10][74]=0;ram[10][75]=0;ram[10][76]=1;ram[10][77]=0;ram[10][78]=0;ram[10][79]=0;ram[10][80]=1;ram[10][81]=0;ram[10][82]=0;ram[10][83]=0;ram[10][84]=0;ram[10][85]=0;ram[10][86]=0;ram[10][87]=0;ram[10][88]=0;ram[10][89]=0;ram[10][90]=0;ram[10][91]=0;ram[10][92]=0;ram[10][93]=0;ram[10][94]=0;ram[10][95]=0;ram[10][96]=0;ram[10][97]=0;ram[10][98]=0;ram[10][99]=0;ram[10][100]=0;ram[10][101]=0;ram[10][102]=0;ram[10][103]=0;ram[10][104]=0;ram[10][105]=0;ram[10][106]=0;ram[10][107]=0;ram[10][108]=0;ram[10][109]=0;ram[10][110]=0;ram[10][111]=0;ram[10][112]=0;ram[10][113]=0;ram[10][114]=0;ram[10][115]=0;ram[10][116]=0;ram[10][117]=0;ram[10][118]=0;ram[10][119]=0;ram[10][120]=0;ram[10][121]=0;ram[10][122]=0;ram[10][123]=0;ram[10][124]=0;ram[10][125]=0;ram[10][126]=0;ram[10][127]=0;ram[10][128]=0;ram[10][129]=0;ram[10][130]=0;ram[10][131]=0;ram[10][132]=0;ram[10][133]=0;ram[10][134]=0;ram[10][135]=0;ram[10][136]=0;ram[10][137]=0;ram[10][138]=0;ram[10][139]=0;ram[10][140]=0;
        ram[11][0]=0;ram[11][1]=0;ram[11][2]=0;ram[11][3]=0;ram[11][4]=0;ram[11][5]=0;ram[11][6]=0;ram[11][7]=0;ram[11][8]=0;ram[11][9]=0;ram[11][10]=0;ram[11][11]=0;ram[11][12]=0;ram[11][13]=0;ram[11][14]=0;ram[11][15]=0;ram[11][16]=0;ram[11][17]=0;ram[11][18]=0;ram[11][19]=0;ram[11][20]=0;ram[11][21]=0;ram[11][22]=0;ram[11][23]=0;ram[11][24]=0;ram[11][25]=0;ram[11][26]=0;ram[11][27]=0;ram[11][28]=0;ram[11][29]=0;ram[11][30]=0;ram[11][31]=0;ram[11][32]=0;ram[11][33]=0;ram[11][34]=0;ram[11][35]=0;ram[11][36]=0;ram[11][37]=0;ram[11][38]=0;ram[11][39]=0;ram[11][40]=0;ram[11][41]=0;ram[11][42]=0;ram[11][43]=0;ram[11][44]=0;ram[11][45]=0;ram[11][46]=0;ram[11][47]=0;ram[11][48]=0;ram[11][49]=0;ram[11][50]=0;ram[11][51]=0;ram[11][52]=0;ram[11][53]=0;ram[11][54]=0;ram[11][55]=0;ram[11][56]=0;ram[11][57]=0;ram[11][58]=0;ram[11][59]=1;ram[11][60]=0;ram[11][61]=1;ram[11][62]=0;ram[11][63]=1;ram[11][64]=0;ram[11][65]=0;ram[11][66]=0;ram[11][67]=0;ram[11][68]=0;ram[11][69]=1;ram[11][70]=0;ram[11][71]=1;ram[11][72]=0;ram[11][73]=1;ram[11][74]=0;ram[11][75]=1;ram[11][76]=0;ram[11][77]=1;ram[11][78]=0;ram[11][79]=1;ram[11][80]=0;ram[11][81]=1;ram[11][82]=0;ram[11][83]=0;ram[11][84]=0;ram[11][85]=0;ram[11][86]=0;ram[11][87]=0;ram[11][88]=0;ram[11][89]=0;ram[11][90]=0;ram[11][91]=0;ram[11][92]=0;ram[11][93]=0;ram[11][94]=0;ram[11][95]=0;ram[11][96]=0;ram[11][97]=0;ram[11][98]=0;ram[11][99]=0;ram[11][100]=0;ram[11][101]=0;ram[11][102]=0;ram[11][103]=0;ram[11][104]=0;ram[11][105]=0;ram[11][106]=0;ram[11][107]=0;ram[11][108]=0;ram[11][109]=0;ram[11][110]=0;ram[11][111]=0;ram[11][112]=0;ram[11][113]=0;ram[11][114]=0;ram[11][115]=0;ram[11][116]=0;ram[11][117]=0;ram[11][118]=0;ram[11][119]=0;ram[11][120]=0;ram[11][121]=0;ram[11][122]=0;ram[11][123]=0;ram[11][124]=0;ram[11][125]=0;ram[11][126]=0;ram[11][127]=0;ram[11][128]=0;ram[11][129]=0;ram[11][130]=0;ram[11][131]=0;ram[11][132]=0;ram[11][133]=0;ram[11][134]=0;ram[11][135]=0;ram[11][136]=0;ram[11][137]=0;ram[11][138]=0;ram[11][139]=0;ram[11][140]=0;
        ram[12][0]=0;ram[12][1]=0;ram[12][2]=0;ram[12][3]=0;ram[12][4]=0;ram[12][5]=0;ram[12][6]=0;ram[12][7]=0;ram[12][8]=0;ram[12][9]=0;ram[12][10]=0;ram[12][11]=0;ram[12][12]=0;ram[12][13]=0;ram[12][14]=0;ram[12][15]=0;ram[12][16]=0;ram[12][17]=0;ram[12][18]=0;ram[12][19]=0;ram[12][20]=0;ram[12][21]=0;ram[12][22]=0;ram[12][23]=0;ram[12][24]=0;ram[12][25]=0;ram[12][26]=0;ram[12][27]=0;ram[12][28]=0;ram[12][29]=0;ram[12][30]=0;ram[12][31]=0;ram[12][32]=0;ram[12][33]=0;ram[12][34]=0;ram[12][35]=0;ram[12][36]=0;ram[12][37]=0;ram[12][38]=0;ram[12][39]=0;ram[12][40]=0;ram[12][41]=0;ram[12][42]=0;ram[12][43]=0;ram[12][44]=0;ram[12][45]=0;ram[12][46]=0;ram[12][47]=0;ram[12][48]=0;ram[12][49]=0;ram[12][50]=0;ram[12][51]=0;ram[12][52]=0;ram[12][53]=0;ram[12][54]=0;ram[12][55]=0;ram[12][56]=0;ram[12][57]=0;ram[12][58]=1;ram[12][59]=0;ram[12][60]=1;ram[12][61]=0;ram[12][62]=1;ram[12][63]=0;ram[12][64]=1;ram[12][65]=0;ram[12][66]=1;ram[12][67]=0;ram[12][68]=1;ram[12][69]=0;ram[12][70]=1;ram[12][71]=0;ram[12][72]=0;ram[12][73]=0;ram[12][74]=0;ram[12][75]=0;ram[12][76]=0;ram[12][77]=0;ram[12][78]=1;ram[12][79]=0;ram[12][80]=1;ram[12][81]=0;ram[12][82]=1;ram[12][83]=0;ram[12][84]=0;ram[12][85]=0;ram[12][86]=0;ram[12][87]=0;ram[12][88]=0;ram[12][89]=0;ram[12][90]=0;ram[12][91]=0;ram[12][92]=0;ram[12][93]=0;ram[12][94]=0;ram[12][95]=0;ram[12][96]=0;ram[12][97]=0;ram[12][98]=0;ram[12][99]=0;ram[12][100]=0;ram[12][101]=0;ram[12][102]=0;ram[12][103]=0;ram[12][104]=0;ram[12][105]=0;ram[12][106]=0;ram[12][107]=0;ram[12][108]=0;ram[12][109]=0;ram[12][110]=0;ram[12][111]=0;ram[12][112]=0;ram[12][113]=0;ram[12][114]=0;ram[12][115]=0;ram[12][116]=0;ram[12][117]=0;ram[12][118]=0;ram[12][119]=0;ram[12][120]=0;ram[12][121]=0;ram[12][122]=0;ram[12][123]=0;ram[12][124]=0;ram[12][125]=0;ram[12][126]=0;ram[12][127]=0;ram[12][128]=0;ram[12][129]=0;ram[12][130]=0;ram[12][131]=0;ram[12][132]=0;ram[12][133]=0;ram[12][134]=0;ram[12][135]=0;ram[12][136]=0;ram[12][137]=0;ram[12][138]=0;ram[12][139]=0;ram[12][140]=0;
        ram[13][0]=0;ram[13][1]=0;ram[13][2]=0;ram[13][3]=0;ram[13][4]=0;ram[13][5]=0;ram[13][6]=0;ram[13][7]=0;ram[13][8]=0;ram[13][9]=0;ram[13][10]=0;ram[13][11]=0;ram[13][12]=0;ram[13][13]=0;ram[13][14]=0;ram[13][15]=0;ram[13][16]=0;ram[13][17]=0;ram[13][18]=0;ram[13][19]=0;ram[13][20]=0;ram[13][21]=0;ram[13][22]=0;ram[13][23]=0;ram[13][24]=0;ram[13][25]=0;ram[13][26]=0;ram[13][27]=0;ram[13][28]=0;ram[13][29]=0;ram[13][30]=0;ram[13][31]=0;ram[13][32]=0;ram[13][33]=0;ram[13][34]=0;ram[13][35]=0;ram[13][36]=0;ram[13][37]=0;ram[13][38]=0;ram[13][39]=0;ram[13][40]=0;ram[13][41]=0;ram[13][42]=0;ram[13][43]=0;ram[13][44]=0;ram[13][45]=0;ram[13][46]=0;ram[13][47]=0;ram[13][48]=0;ram[13][49]=0;ram[13][50]=0;ram[13][51]=0;ram[13][52]=0;ram[13][53]=0;ram[13][54]=0;ram[13][55]=0;ram[13][56]=0;ram[13][57]=1;ram[13][58]=0;ram[13][59]=1;ram[13][60]=0;ram[13][61]=1;ram[13][62]=0;ram[13][63]=0;ram[13][64]=0;ram[13][65]=1;ram[13][66]=0;ram[13][67]=1;ram[13][68]=0;ram[13][69]=1;ram[13][70]=0;ram[13][71]=0;ram[13][72]=0;ram[13][73]=1;ram[13][74]=0;ram[13][75]=1;ram[13][76]=0;ram[13][77]=1;ram[13][78]=0;ram[13][79]=1;ram[13][80]=0;ram[13][81]=0;ram[13][82]=0;ram[13][83]=1;ram[13][84]=0;ram[13][85]=0;ram[13][86]=0;ram[13][87]=0;ram[13][88]=0;ram[13][89]=0;ram[13][90]=0;ram[13][91]=0;ram[13][92]=0;ram[13][93]=0;ram[13][94]=0;ram[13][95]=0;ram[13][96]=0;ram[13][97]=0;ram[13][98]=0;ram[13][99]=0;ram[13][100]=0;ram[13][101]=0;ram[13][102]=0;ram[13][103]=0;ram[13][104]=0;ram[13][105]=0;ram[13][106]=0;ram[13][107]=0;ram[13][108]=0;ram[13][109]=0;ram[13][110]=0;ram[13][111]=0;ram[13][112]=0;ram[13][113]=0;ram[13][114]=0;ram[13][115]=0;ram[13][116]=0;ram[13][117]=0;ram[13][118]=0;ram[13][119]=0;ram[13][120]=0;ram[13][121]=0;ram[13][122]=0;ram[13][123]=0;ram[13][124]=0;ram[13][125]=0;ram[13][126]=0;ram[13][127]=0;ram[13][128]=0;ram[13][129]=0;ram[13][130]=0;ram[13][131]=0;ram[13][132]=0;ram[13][133]=0;ram[13][134]=0;ram[13][135]=0;ram[13][136]=0;ram[13][137]=0;ram[13][138]=0;ram[13][139]=0;ram[13][140]=0;
        ram[14][0]=0;ram[14][1]=0;ram[14][2]=0;ram[14][3]=0;ram[14][4]=0;ram[14][5]=0;ram[14][6]=0;ram[14][7]=0;ram[14][8]=0;ram[14][9]=0;ram[14][10]=0;ram[14][11]=0;ram[14][12]=0;ram[14][13]=0;ram[14][14]=0;ram[14][15]=0;ram[14][16]=0;ram[14][17]=0;ram[14][18]=0;ram[14][19]=0;ram[14][20]=0;ram[14][21]=0;ram[14][22]=0;ram[14][23]=0;ram[14][24]=0;ram[14][25]=0;ram[14][26]=0;ram[14][27]=0;ram[14][28]=0;ram[14][29]=0;ram[14][30]=0;ram[14][31]=0;ram[14][32]=0;ram[14][33]=0;ram[14][34]=0;ram[14][35]=0;ram[14][36]=0;ram[14][37]=0;ram[14][38]=0;ram[14][39]=0;ram[14][40]=0;ram[14][41]=0;ram[14][42]=0;ram[14][43]=0;ram[14][44]=0;ram[14][45]=0;ram[14][46]=0;ram[14][47]=0;ram[14][48]=0;ram[14][49]=0;ram[14][50]=0;ram[14][51]=0;ram[14][52]=0;ram[14][53]=0;ram[14][54]=0;ram[14][55]=0;ram[14][56]=1;ram[14][57]=0;ram[14][58]=1;ram[14][59]=0;ram[14][60]=1;ram[14][61]=0;ram[14][62]=0;ram[14][63]=0;ram[14][64]=1;ram[14][65]=0;ram[14][66]=0;ram[14][67]=0;ram[14][68]=1;ram[14][69]=0;ram[14][70]=1;ram[14][71]=0;ram[14][72]=1;ram[14][73]=0;ram[14][74]=1;ram[14][75]=0;ram[14][76]=1;ram[14][77]=0;ram[14][78]=1;ram[14][79]=0;ram[14][80]=1;ram[14][81]=0;ram[14][82]=1;ram[14][83]=0;ram[14][84]=1;ram[14][85]=0;ram[14][86]=0;ram[14][87]=0;ram[14][88]=0;ram[14][89]=0;ram[14][90]=0;ram[14][91]=0;ram[14][92]=0;ram[14][93]=0;ram[14][94]=0;ram[14][95]=0;ram[14][96]=0;ram[14][97]=0;ram[14][98]=0;ram[14][99]=0;ram[14][100]=0;ram[14][101]=0;ram[14][102]=0;ram[14][103]=0;ram[14][104]=0;ram[14][105]=0;ram[14][106]=0;ram[14][107]=0;ram[14][108]=0;ram[14][109]=0;ram[14][110]=0;ram[14][111]=0;ram[14][112]=0;ram[14][113]=0;ram[14][114]=0;ram[14][115]=0;ram[14][116]=0;ram[14][117]=0;ram[14][118]=0;ram[14][119]=0;ram[14][120]=0;ram[14][121]=0;ram[14][122]=0;ram[14][123]=0;ram[14][124]=0;ram[14][125]=0;ram[14][126]=0;ram[14][127]=0;ram[14][128]=0;ram[14][129]=0;ram[14][130]=0;ram[14][131]=0;ram[14][132]=0;ram[14][133]=0;ram[14][134]=0;ram[14][135]=0;ram[14][136]=0;ram[14][137]=0;ram[14][138]=0;ram[14][139]=0;ram[14][140]=0;
        ram[15][0]=0;ram[15][1]=0;ram[15][2]=0;ram[15][3]=0;ram[15][4]=0;ram[15][5]=0;ram[15][6]=0;ram[15][7]=0;ram[15][8]=0;ram[15][9]=0;ram[15][10]=0;ram[15][11]=0;ram[15][12]=0;ram[15][13]=0;ram[15][14]=0;ram[15][15]=0;ram[15][16]=0;ram[15][17]=0;ram[15][18]=0;ram[15][19]=0;ram[15][20]=0;ram[15][21]=0;ram[15][22]=0;ram[15][23]=0;ram[15][24]=0;ram[15][25]=0;ram[15][26]=0;ram[15][27]=0;ram[15][28]=0;ram[15][29]=0;ram[15][30]=0;ram[15][31]=0;ram[15][32]=0;ram[15][33]=0;ram[15][34]=0;ram[15][35]=0;ram[15][36]=0;ram[15][37]=0;ram[15][38]=0;ram[15][39]=0;ram[15][40]=0;ram[15][41]=0;ram[15][42]=0;ram[15][43]=0;ram[15][44]=0;ram[15][45]=0;ram[15][46]=0;ram[15][47]=0;ram[15][48]=0;ram[15][49]=0;ram[15][50]=0;ram[15][51]=0;ram[15][52]=0;ram[15][53]=0;ram[15][54]=0;ram[15][55]=1;ram[15][56]=0;ram[15][57]=1;ram[15][58]=0;ram[15][59]=0;ram[15][60]=0;ram[15][61]=1;ram[15][62]=0;ram[15][63]=1;ram[15][64]=0;ram[15][65]=1;ram[15][66]=0;ram[15][67]=1;ram[15][68]=0;ram[15][69]=1;ram[15][70]=0;ram[15][71]=0;ram[15][72]=0;ram[15][73]=1;ram[15][74]=0;ram[15][75]=1;ram[15][76]=0;ram[15][77]=1;ram[15][78]=0;ram[15][79]=1;ram[15][80]=0;ram[15][81]=0;ram[15][82]=0;ram[15][83]=0;ram[15][84]=0;ram[15][85]=1;ram[15][86]=0;ram[15][87]=0;ram[15][88]=0;ram[15][89]=0;ram[15][90]=0;ram[15][91]=0;ram[15][92]=0;ram[15][93]=0;ram[15][94]=0;ram[15][95]=0;ram[15][96]=0;ram[15][97]=0;ram[15][98]=0;ram[15][99]=0;ram[15][100]=0;ram[15][101]=0;ram[15][102]=0;ram[15][103]=0;ram[15][104]=0;ram[15][105]=0;ram[15][106]=0;ram[15][107]=0;ram[15][108]=0;ram[15][109]=0;ram[15][110]=0;ram[15][111]=0;ram[15][112]=0;ram[15][113]=0;ram[15][114]=0;ram[15][115]=0;ram[15][116]=0;ram[15][117]=0;ram[15][118]=0;ram[15][119]=0;ram[15][120]=0;ram[15][121]=0;ram[15][122]=0;ram[15][123]=0;ram[15][124]=0;ram[15][125]=0;ram[15][126]=0;ram[15][127]=0;ram[15][128]=0;ram[15][129]=0;ram[15][130]=0;ram[15][131]=0;ram[15][132]=0;ram[15][133]=0;ram[15][134]=0;ram[15][135]=0;ram[15][136]=0;ram[15][137]=0;ram[15][138]=0;ram[15][139]=0;ram[15][140]=0;
        ram[16][0]=0;ram[16][1]=0;ram[16][2]=0;ram[16][3]=0;ram[16][4]=0;ram[16][5]=0;ram[16][6]=0;ram[16][7]=0;ram[16][8]=0;ram[16][9]=0;ram[16][10]=0;ram[16][11]=0;ram[16][12]=0;ram[16][13]=0;ram[16][14]=0;ram[16][15]=0;ram[16][16]=0;ram[16][17]=0;ram[16][18]=0;ram[16][19]=0;ram[16][20]=0;ram[16][21]=0;ram[16][22]=0;ram[16][23]=0;ram[16][24]=0;ram[16][25]=0;ram[16][26]=0;ram[16][27]=0;ram[16][28]=0;ram[16][29]=0;ram[16][30]=0;ram[16][31]=0;ram[16][32]=0;ram[16][33]=0;ram[16][34]=0;ram[16][35]=0;ram[16][36]=0;ram[16][37]=0;ram[16][38]=0;ram[16][39]=0;ram[16][40]=0;ram[16][41]=0;ram[16][42]=0;ram[16][43]=0;ram[16][44]=0;ram[16][45]=0;ram[16][46]=0;ram[16][47]=0;ram[16][48]=0;ram[16][49]=0;ram[16][50]=0;ram[16][51]=0;ram[16][52]=0;ram[16][53]=0;ram[16][54]=1;ram[16][55]=0;ram[16][56]=0;ram[16][57]=0;ram[16][58]=1;ram[16][59]=0;ram[16][60]=1;ram[16][61]=0;ram[16][62]=0;ram[16][63]=0;ram[16][64]=1;ram[16][65]=0;ram[16][66]=1;ram[16][67]=0;ram[16][68]=1;ram[16][69]=0;ram[16][70]=1;ram[16][71]=0;ram[16][72]=1;ram[16][73]=0;ram[16][74]=1;ram[16][75]=0;ram[16][76]=0;ram[16][77]=0;ram[16][78]=1;ram[16][79]=0;ram[16][80]=0;ram[16][81]=0;ram[16][82]=1;ram[16][83]=0;ram[16][84]=1;ram[16][85]=0;ram[16][86]=1;ram[16][87]=0;ram[16][88]=0;ram[16][89]=0;ram[16][90]=0;ram[16][91]=0;ram[16][92]=0;ram[16][93]=0;ram[16][94]=0;ram[16][95]=0;ram[16][96]=0;ram[16][97]=0;ram[16][98]=0;ram[16][99]=0;ram[16][100]=0;ram[16][101]=0;ram[16][102]=0;ram[16][103]=0;ram[16][104]=0;ram[16][105]=0;ram[16][106]=0;ram[16][107]=0;ram[16][108]=0;ram[16][109]=0;ram[16][110]=0;ram[16][111]=0;ram[16][112]=0;ram[16][113]=0;ram[16][114]=0;ram[16][115]=0;ram[16][116]=0;ram[16][117]=0;ram[16][118]=0;ram[16][119]=0;ram[16][120]=0;ram[16][121]=0;ram[16][122]=0;ram[16][123]=0;ram[16][124]=0;ram[16][125]=0;ram[16][126]=0;ram[16][127]=0;ram[16][128]=0;ram[16][129]=0;ram[16][130]=0;ram[16][131]=0;ram[16][132]=0;ram[16][133]=0;ram[16][134]=0;ram[16][135]=0;ram[16][136]=0;ram[16][137]=0;ram[16][138]=0;ram[16][139]=0;ram[16][140]=0;
        ram[17][0]=0;ram[17][1]=0;ram[17][2]=0;ram[17][3]=0;ram[17][4]=0;ram[17][5]=0;ram[17][6]=0;ram[17][7]=0;ram[17][8]=0;ram[17][9]=0;ram[17][10]=0;ram[17][11]=0;ram[17][12]=0;ram[17][13]=0;ram[17][14]=0;ram[17][15]=0;ram[17][16]=0;ram[17][17]=0;ram[17][18]=0;ram[17][19]=0;ram[17][20]=0;ram[17][21]=0;ram[17][22]=0;ram[17][23]=0;ram[17][24]=0;ram[17][25]=0;ram[17][26]=0;ram[17][27]=0;ram[17][28]=0;ram[17][29]=0;ram[17][30]=0;ram[17][31]=0;ram[17][32]=0;ram[17][33]=0;ram[17][34]=0;ram[17][35]=0;ram[17][36]=0;ram[17][37]=0;ram[17][38]=0;ram[17][39]=0;ram[17][40]=0;ram[17][41]=0;ram[17][42]=0;ram[17][43]=0;ram[17][44]=0;ram[17][45]=0;ram[17][46]=0;ram[17][47]=0;ram[17][48]=0;ram[17][49]=0;ram[17][50]=0;ram[17][51]=0;ram[17][52]=0;ram[17][53]=1;ram[17][54]=0;ram[17][55]=1;ram[17][56]=0;ram[17][57]=1;ram[17][58]=0;ram[17][59]=1;ram[17][60]=0;ram[17][61]=0;ram[17][62]=0;ram[17][63]=1;ram[17][64]=0;ram[17][65]=0;ram[17][66]=0;ram[17][67]=1;ram[17][68]=0;ram[17][69]=1;ram[17][70]=0;ram[17][71]=1;ram[17][72]=0;ram[17][73]=1;ram[17][74]=0;ram[17][75]=1;ram[17][76]=0;ram[17][77]=1;ram[17][78]=0;ram[17][79]=1;ram[17][80]=0;ram[17][81]=1;ram[17][82]=0;ram[17][83]=0;ram[17][84]=0;ram[17][85]=0;ram[17][86]=0;ram[17][87]=1;ram[17][88]=0;ram[17][89]=0;ram[17][90]=0;ram[17][91]=0;ram[17][92]=0;ram[17][93]=0;ram[17][94]=0;ram[17][95]=0;ram[17][96]=0;ram[17][97]=0;ram[17][98]=0;ram[17][99]=0;ram[17][100]=0;ram[17][101]=0;ram[17][102]=0;ram[17][103]=0;ram[17][104]=0;ram[17][105]=0;ram[17][106]=0;ram[17][107]=0;ram[17][108]=0;ram[17][109]=0;ram[17][110]=0;ram[17][111]=0;ram[17][112]=0;ram[17][113]=0;ram[17][114]=0;ram[17][115]=0;ram[17][116]=0;ram[17][117]=0;ram[17][118]=0;ram[17][119]=0;ram[17][120]=0;ram[17][121]=0;ram[17][122]=0;ram[17][123]=0;ram[17][124]=0;ram[17][125]=0;ram[17][126]=0;ram[17][127]=0;ram[17][128]=0;ram[17][129]=0;ram[17][130]=0;ram[17][131]=0;ram[17][132]=0;ram[17][133]=0;ram[17][134]=0;ram[17][135]=0;ram[17][136]=0;ram[17][137]=0;ram[17][138]=0;ram[17][139]=0;ram[17][140]=0;
        ram[18][0]=0;ram[18][1]=0;ram[18][2]=0;ram[18][3]=0;ram[18][4]=0;ram[18][5]=0;ram[18][6]=0;ram[18][7]=0;ram[18][8]=0;ram[18][9]=0;ram[18][10]=0;ram[18][11]=0;ram[18][12]=0;ram[18][13]=0;ram[18][14]=0;ram[18][15]=0;ram[18][16]=0;ram[18][17]=0;ram[18][18]=0;ram[18][19]=0;ram[18][20]=0;ram[18][21]=0;ram[18][22]=0;ram[18][23]=0;ram[18][24]=0;ram[18][25]=0;ram[18][26]=0;ram[18][27]=0;ram[18][28]=0;ram[18][29]=0;ram[18][30]=0;ram[18][31]=0;ram[18][32]=0;ram[18][33]=0;ram[18][34]=0;ram[18][35]=0;ram[18][36]=0;ram[18][37]=0;ram[18][38]=0;ram[18][39]=0;ram[18][40]=0;ram[18][41]=0;ram[18][42]=0;ram[18][43]=0;ram[18][44]=0;ram[18][45]=0;ram[18][46]=0;ram[18][47]=0;ram[18][48]=0;ram[18][49]=0;ram[18][50]=0;ram[18][51]=0;ram[18][52]=1;ram[18][53]=0;ram[18][54]=0;ram[18][55]=0;ram[18][56]=0;ram[18][57]=0;ram[18][58]=1;ram[18][59]=0;ram[18][60]=1;ram[18][61]=0;ram[18][62]=0;ram[18][63]=0;ram[18][64]=0;ram[18][65]=0;ram[18][66]=1;ram[18][67]=0;ram[18][68]=1;ram[18][69]=0;ram[18][70]=0;ram[18][71]=0;ram[18][72]=1;ram[18][73]=0;ram[18][74]=1;ram[18][75]=0;ram[18][76]=1;ram[18][77]=0;ram[18][78]=0;ram[18][79]=0;ram[18][80]=1;ram[18][81]=0;ram[18][82]=1;ram[18][83]=0;ram[18][84]=0;ram[18][85]=0;ram[18][86]=1;ram[18][87]=0;ram[18][88]=1;ram[18][89]=0;ram[18][90]=0;ram[18][91]=0;ram[18][92]=0;ram[18][93]=0;ram[18][94]=0;ram[18][95]=0;ram[18][96]=0;ram[18][97]=0;ram[18][98]=0;ram[18][99]=0;ram[18][100]=0;ram[18][101]=0;ram[18][102]=0;ram[18][103]=0;ram[18][104]=0;ram[18][105]=0;ram[18][106]=0;ram[18][107]=0;ram[18][108]=0;ram[18][109]=0;ram[18][110]=0;ram[18][111]=0;ram[18][112]=0;ram[18][113]=0;ram[18][114]=0;ram[18][115]=0;ram[18][116]=0;ram[18][117]=0;ram[18][118]=0;ram[18][119]=0;ram[18][120]=0;ram[18][121]=0;ram[18][122]=0;ram[18][123]=0;ram[18][124]=0;ram[18][125]=0;ram[18][126]=0;ram[18][127]=0;ram[18][128]=0;ram[18][129]=0;ram[18][130]=0;ram[18][131]=0;ram[18][132]=0;ram[18][133]=0;ram[18][134]=0;ram[18][135]=0;ram[18][136]=0;ram[18][137]=0;ram[18][138]=0;ram[18][139]=0;ram[18][140]=0;
        ram[19][0]=0;ram[19][1]=0;ram[19][2]=0;ram[19][3]=0;ram[19][4]=0;ram[19][5]=0;ram[19][6]=0;ram[19][7]=0;ram[19][8]=0;ram[19][9]=0;ram[19][10]=0;ram[19][11]=0;ram[19][12]=0;ram[19][13]=0;ram[19][14]=0;ram[19][15]=0;ram[19][16]=0;ram[19][17]=0;ram[19][18]=0;ram[19][19]=0;ram[19][20]=0;ram[19][21]=0;ram[19][22]=0;ram[19][23]=0;ram[19][24]=0;ram[19][25]=0;ram[19][26]=0;ram[19][27]=0;ram[19][28]=0;ram[19][29]=0;ram[19][30]=0;ram[19][31]=0;ram[19][32]=0;ram[19][33]=0;ram[19][34]=0;ram[19][35]=0;ram[19][36]=0;ram[19][37]=0;ram[19][38]=0;ram[19][39]=0;ram[19][40]=0;ram[19][41]=0;ram[19][42]=0;ram[19][43]=0;ram[19][44]=0;ram[19][45]=0;ram[19][46]=0;ram[19][47]=0;ram[19][48]=0;ram[19][49]=0;ram[19][50]=0;ram[19][51]=1;ram[19][52]=0;ram[19][53]=0;ram[19][54]=0;ram[19][55]=1;ram[19][56]=0;ram[19][57]=0;ram[19][58]=0;ram[19][59]=0;ram[19][60]=0;ram[19][61]=1;ram[19][62]=0;ram[19][63]=1;ram[19][64]=0;ram[19][65]=0;ram[19][66]=0;ram[19][67]=1;ram[19][68]=0;ram[19][69]=1;ram[19][70]=0;ram[19][71]=1;ram[19][72]=0;ram[19][73]=1;ram[19][74]=0;ram[19][75]=0;ram[19][76]=0;ram[19][77]=1;ram[19][78]=0;ram[19][79]=1;ram[19][80]=0;ram[19][81]=1;ram[19][82]=0;ram[19][83]=1;ram[19][84]=0;ram[19][85]=0;ram[19][86]=0;ram[19][87]=1;ram[19][88]=0;ram[19][89]=1;ram[19][90]=0;ram[19][91]=0;ram[19][92]=0;ram[19][93]=0;ram[19][94]=0;ram[19][95]=0;ram[19][96]=0;ram[19][97]=0;ram[19][98]=0;ram[19][99]=0;ram[19][100]=0;ram[19][101]=0;ram[19][102]=0;ram[19][103]=0;ram[19][104]=0;ram[19][105]=0;ram[19][106]=0;ram[19][107]=0;ram[19][108]=0;ram[19][109]=0;ram[19][110]=0;ram[19][111]=0;ram[19][112]=0;ram[19][113]=0;ram[19][114]=0;ram[19][115]=0;ram[19][116]=0;ram[19][117]=0;ram[19][118]=0;ram[19][119]=0;ram[19][120]=0;ram[19][121]=0;ram[19][122]=0;ram[19][123]=0;ram[19][124]=0;ram[19][125]=0;ram[19][126]=0;ram[19][127]=0;ram[19][128]=0;ram[19][129]=0;ram[19][130]=0;ram[19][131]=0;ram[19][132]=0;ram[19][133]=0;ram[19][134]=0;ram[19][135]=0;ram[19][136]=0;ram[19][137]=0;ram[19][138]=0;ram[19][139]=0;ram[19][140]=0;
        ram[20][0]=0;ram[20][1]=0;ram[20][2]=0;ram[20][3]=0;ram[20][4]=0;ram[20][5]=0;ram[20][6]=0;ram[20][7]=0;ram[20][8]=0;ram[20][9]=0;ram[20][10]=0;ram[20][11]=0;ram[20][12]=0;ram[20][13]=0;ram[20][14]=0;ram[20][15]=0;ram[20][16]=0;ram[20][17]=0;ram[20][18]=0;ram[20][19]=0;ram[20][20]=0;ram[20][21]=0;ram[20][22]=0;ram[20][23]=0;ram[20][24]=0;ram[20][25]=0;ram[20][26]=0;ram[20][27]=0;ram[20][28]=0;ram[20][29]=0;ram[20][30]=0;ram[20][31]=0;ram[20][32]=0;ram[20][33]=0;ram[20][34]=0;ram[20][35]=0;ram[20][36]=0;ram[20][37]=0;ram[20][38]=0;ram[20][39]=0;ram[20][40]=0;ram[20][41]=0;ram[20][42]=0;ram[20][43]=0;ram[20][44]=0;ram[20][45]=0;ram[20][46]=0;ram[20][47]=0;ram[20][48]=0;ram[20][49]=0;ram[20][50]=1;ram[20][51]=0;ram[20][52]=1;ram[20][53]=0;ram[20][54]=1;ram[20][55]=0;ram[20][56]=1;ram[20][57]=0;ram[20][58]=0;ram[20][59]=0;ram[20][60]=1;ram[20][61]=0;ram[20][62]=0;ram[20][63]=0;ram[20][64]=0;ram[20][65]=0;ram[20][66]=0;ram[20][67]=0;ram[20][68]=1;ram[20][69]=0;ram[20][70]=0;ram[20][71]=0;ram[20][72]=0;ram[20][73]=0;ram[20][74]=1;ram[20][75]=0;ram[20][76]=1;ram[20][77]=0;ram[20][78]=1;ram[20][79]=0;ram[20][80]=0;ram[20][81]=0;ram[20][82]=0;ram[20][83]=0;ram[20][84]=1;ram[20][85]=0;ram[20][86]=0;ram[20][87]=0;ram[20][88]=1;ram[20][89]=0;ram[20][90]=1;ram[20][91]=0;ram[20][92]=0;ram[20][93]=0;ram[20][94]=0;ram[20][95]=0;ram[20][96]=0;ram[20][97]=0;ram[20][98]=0;ram[20][99]=0;ram[20][100]=0;ram[20][101]=0;ram[20][102]=0;ram[20][103]=0;ram[20][104]=0;ram[20][105]=0;ram[20][106]=0;ram[20][107]=0;ram[20][108]=0;ram[20][109]=0;ram[20][110]=0;ram[20][111]=0;ram[20][112]=0;ram[20][113]=0;ram[20][114]=0;ram[20][115]=0;ram[20][116]=0;ram[20][117]=0;ram[20][118]=0;ram[20][119]=0;ram[20][120]=0;ram[20][121]=0;ram[20][122]=0;ram[20][123]=0;ram[20][124]=0;ram[20][125]=0;ram[20][126]=0;ram[20][127]=0;ram[20][128]=0;ram[20][129]=0;ram[20][130]=0;ram[20][131]=0;ram[20][132]=0;ram[20][133]=0;ram[20][134]=0;ram[20][135]=0;ram[20][136]=0;ram[20][137]=0;ram[20][138]=0;ram[20][139]=0;ram[20][140]=0;
        ram[21][0]=0;ram[21][1]=0;ram[21][2]=0;ram[21][3]=0;ram[21][4]=0;ram[21][5]=0;ram[21][6]=0;ram[21][7]=0;ram[21][8]=0;ram[21][9]=0;ram[21][10]=0;ram[21][11]=0;ram[21][12]=0;ram[21][13]=0;ram[21][14]=0;ram[21][15]=0;ram[21][16]=0;ram[21][17]=0;ram[21][18]=0;ram[21][19]=0;ram[21][20]=0;ram[21][21]=0;ram[21][22]=0;ram[21][23]=0;ram[21][24]=0;ram[21][25]=0;ram[21][26]=0;ram[21][27]=0;ram[21][28]=0;ram[21][29]=0;ram[21][30]=0;ram[21][31]=0;ram[21][32]=0;ram[21][33]=0;ram[21][34]=0;ram[21][35]=0;ram[21][36]=0;ram[21][37]=0;ram[21][38]=0;ram[21][39]=0;ram[21][40]=0;ram[21][41]=0;ram[21][42]=0;ram[21][43]=0;ram[21][44]=0;ram[21][45]=0;ram[21][46]=0;ram[21][47]=0;ram[21][48]=0;ram[21][49]=1;ram[21][50]=0;ram[21][51]=1;ram[21][52]=0;ram[21][53]=1;ram[21][54]=0;ram[21][55]=0;ram[21][56]=0;ram[21][57]=0;ram[21][58]=0;ram[21][59]=1;ram[21][60]=0;ram[21][61]=1;ram[21][62]=0;ram[21][63]=1;ram[21][64]=0;ram[21][65]=1;ram[21][66]=0;ram[21][67]=1;ram[21][68]=0;ram[21][69]=1;ram[21][70]=0;ram[21][71]=1;ram[21][72]=0;ram[21][73]=1;ram[21][74]=0;ram[21][75]=1;ram[21][76]=0;ram[21][77]=1;ram[21][78]=0;ram[21][79]=1;ram[21][80]=0;ram[21][81]=1;ram[21][82]=0;ram[21][83]=1;ram[21][84]=0;ram[21][85]=1;ram[21][86]=0;ram[21][87]=0;ram[21][88]=0;ram[21][89]=1;ram[21][90]=0;ram[21][91]=1;ram[21][92]=0;ram[21][93]=0;ram[21][94]=0;ram[21][95]=0;ram[21][96]=0;ram[21][97]=0;ram[21][98]=0;ram[21][99]=0;ram[21][100]=0;ram[21][101]=0;ram[21][102]=0;ram[21][103]=0;ram[21][104]=0;ram[21][105]=0;ram[21][106]=0;ram[21][107]=0;ram[21][108]=0;ram[21][109]=0;ram[21][110]=0;ram[21][111]=0;ram[21][112]=0;ram[21][113]=0;ram[21][114]=0;ram[21][115]=0;ram[21][116]=0;ram[21][117]=0;ram[21][118]=0;ram[21][119]=0;ram[21][120]=0;ram[21][121]=0;ram[21][122]=0;ram[21][123]=0;ram[21][124]=0;ram[21][125]=0;ram[21][126]=0;ram[21][127]=0;ram[21][128]=0;ram[21][129]=0;ram[21][130]=0;ram[21][131]=0;ram[21][132]=0;ram[21][133]=0;ram[21][134]=0;ram[21][135]=0;ram[21][136]=0;ram[21][137]=0;ram[21][138]=0;ram[21][139]=0;ram[21][140]=0;
        ram[22][0]=0;ram[22][1]=0;ram[22][2]=0;ram[22][3]=0;ram[22][4]=0;ram[22][5]=0;ram[22][6]=0;ram[22][7]=0;ram[22][8]=0;ram[22][9]=0;ram[22][10]=0;ram[22][11]=0;ram[22][12]=0;ram[22][13]=0;ram[22][14]=0;ram[22][15]=0;ram[22][16]=0;ram[22][17]=0;ram[22][18]=0;ram[22][19]=0;ram[22][20]=0;ram[22][21]=0;ram[22][22]=0;ram[22][23]=0;ram[22][24]=0;ram[22][25]=0;ram[22][26]=0;ram[22][27]=0;ram[22][28]=0;ram[22][29]=0;ram[22][30]=0;ram[22][31]=0;ram[22][32]=0;ram[22][33]=0;ram[22][34]=0;ram[22][35]=0;ram[22][36]=0;ram[22][37]=0;ram[22][38]=0;ram[22][39]=0;ram[22][40]=0;ram[22][41]=0;ram[22][42]=0;ram[22][43]=0;ram[22][44]=0;ram[22][45]=0;ram[22][46]=0;ram[22][47]=0;ram[22][48]=1;ram[22][49]=0;ram[22][50]=1;ram[22][51]=0;ram[22][52]=0;ram[22][53]=0;ram[22][54]=1;ram[22][55]=0;ram[22][56]=1;ram[22][57]=0;ram[22][58]=1;ram[22][59]=0;ram[22][60]=0;ram[22][61]=0;ram[22][62]=1;ram[22][63]=0;ram[22][64]=1;ram[22][65]=0;ram[22][66]=0;ram[22][67]=0;ram[22][68]=1;ram[22][69]=0;ram[22][70]=0;ram[22][71]=0;ram[22][72]=1;ram[22][73]=0;ram[22][74]=1;ram[22][75]=0;ram[22][76]=0;ram[22][77]=0;ram[22][78]=1;ram[22][79]=0;ram[22][80]=0;ram[22][81]=0;ram[22][82]=0;ram[22][83]=0;ram[22][84]=1;ram[22][85]=0;ram[22][86]=0;ram[22][87]=0;ram[22][88]=0;ram[22][89]=0;ram[22][90]=1;ram[22][91]=0;ram[22][92]=1;ram[22][93]=0;ram[22][94]=0;ram[22][95]=0;ram[22][96]=0;ram[22][97]=0;ram[22][98]=0;ram[22][99]=0;ram[22][100]=0;ram[22][101]=0;ram[22][102]=0;ram[22][103]=0;ram[22][104]=0;ram[22][105]=0;ram[22][106]=0;ram[22][107]=0;ram[22][108]=0;ram[22][109]=0;ram[22][110]=0;ram[22][111]=0;ram[22][112]=0;ram[22][113]=0;ram[22][114]=0;ram[22][115]=0;ram[22][116]=0;ram[22][117]=0;ram[22][118]=0;ram[22][119]=0;ram[22][120]=0;ram[22][121]=0;ram[22][122]=0;ram[22][123]=0;ram[22][124]=0;ram[22][125]=0;ram[22][126]=0;ram[22][127]=0;ram[22][128]=0;ram[22][129]=0;ram[22][130]=0;ram[22][131]=0;ram[22][132]=0;ram[22][133]=0;ram[22][134]=0;ram[22][135]=0;ram[22][136]=0;ram[22][137]=0;ram[22][138]=0;ram[22][139]=0;ram[22][140]=0;
        ram[23][0]=0;ram[23][1]=0;ram[23][2]=0;ram[23][3]=0;ram[23][4]=0;ram[23][5]=0;ram[23][6]=0;ram[23][7]=0;ram[23][8]=0;ram[23][9]=0;ram[23][10]=0;ram[23][11]=0;ram[23][12]=0;ram[23][13]=0;ram[23][14]=0;ram[23][15]=0;ram[23][16]=0;ram[23][17]=0;ram[23][18]=0;ram[23][19]=0;ram[23][20]=0;ram[23][21]=0;ram[23][22]=0;ram[23][23]=0;ram[23][24]=0;ram[23][25]=0;ram[23][26]=0;ram[23][27]=0;ram[23][28]=0;ram[23][29]=0;ram[23][30]=0;ram[23][31]=0;ram[23][32]=0;ram[23][33]=0;ram[23][34]=0;ram[23][35]=0;ram[23][36]=0;ram[23][37]=0;ram[23][38]=0;ram[23][39]=0;ram[23][40]=0;ram[23][41]=0;ram[23][42]=0;ram[23][43]=0;ram[23][44]=0;ram[23][45]=0;ram[23][46]=0;ram[23][47]=1;ram[23][48]=0;ram[23][49]=1;ram[23][50]=0;ram[23][51]=1;ram[23][52]=0;ram[23][53]=0;ram[23][54]=0;ram[23][55]=1;ram[23][56]=0;ram[23][57]=0;ram[23][58]=0;ram[23][59]=1;ram[23][60]=0;ram[23][61]=1;ram[23][62]=0;ram[23][63]=1;ram[23][64]=0;ram[23][65]=0;ram[23][66]=0;ram[23][67]=0;ram[23][68]=0;ram[23][69]=1;ram[23][70]=0;ram[23][71]=1;ram[23][72]=0;ram[23][73]=1;ram[23][74]=0;ram[23][75]=1;ram[23][76]=0;ram[23][77]=1;ram[23][78]=0;ram[23][79]=1;ram[23][80]=0;ram[23][81]=1;ram[23][82]=0;ram[23][83]=1;ram[23][84]=0;ram[23][85]=1;ram[23][86]=0;ram[23][87]=1;ram[23][88]=0;ram[23][89]=0;ram[23][90]=0;ram[23][91]=0;ram[23][92]=0;ram[23][93]=1;ram[23][94]=0;ram[23][95]=0;ram[23][96]=0;ram[23][97]=0;ram[23][98]=0;ram[23][99]=0;ram[23][100]=0;ram[23][101]=0;ram[23][102]=0;ram[23][103]=0;ram[23][104]=0;ram[23][105]=0;ram[23][106]=0;ram[23][107]=0;ram[23][108]=0;ram[23][109]=0;ram[23][110]=0;ram[23][111]=0;ram[23][112]=0;ram[23][113]=0;ram[23][114]=0;ram[23][115]=0;ram[23][116]=0;ram[23][117]=0;ram[23][118]=0;ram[23][119]=0;ram[23][120]=0;ram[23][121]=0;ram[23][122]=0;ram[23][123]=0;ram[23][124]=0;ram[23][125]=0;ram[23][126]=0;ram[23][127]=0;ram[23][128]=0;ram[23][129]=0;ram[23][130]=0;ram[23][131]=0;ram[23][132]=0;ram[23][133]=0;ram[23][134]=0;ram[23][135]=0;ram[23][136]=0;ram[23][137]=0;ram[23][138]=0;ram[23][139]=0;ram[23][140]=0;
        ram[24][0]=0;ram[24][1]=0;ram[24][2]=0;ram[24][3]=0;ram[24][4]=0;ram[24][5]=0;ram[24][6]=0;ram[24][7]=0;ram[24][8]=0;ram[24][9]=0;ram[24][10]=0;ram[24][11]=0;ram[24][12]=0;ram[24][13]=0;ram[24][14]=0;ram[24][15]=0;ram[24][16]=0;ram[24][17]=0;ram[24][18]=0;ram[24][19]=0;ram[24][20]=0;ram[24][21]=0;ram[24][22]=0;ram[24][23]=0;ram[24][24]=0;ram[24][25]=0;ram[24][26]=0;ram[24][27]=0;ram[24][28]=0;ram[24][29]=0;ram[24][30]=0;ram[24][31]=0;ram[24][32]=0;ram[24][33]=0;ram[24][34]=0;ram[24][35]=0;ram[24][36]=0;ram[24][37]=0;ram[24][38]=0;ram[24][39]=0;ram[24][40]=0;ram[24][41]=0;ram[24][42]=0;ram[24][43]=0;ram[24][44]=0;ram[24][45]=0;ram[24][46]=1;ram[24][47]=0;ram[24][48]=0;ram[24][49]=0;ram[24][50]=1;ram[24][51]=0;ram[24][52]=1;ram[24][53]=0;ram[24][54]=1;ram[24][55]=0;ram[24][56]=1;ram[24][57]=0;ram[24][58]=1;ram[24][59]=0;ram[24][60]=1;ram[24][61]=0;ram[24][62]=1;ram[24][63]=0;ram[24][64]=1;ram[24][65]=0;ram[24][66]=0;ram[24][67]=0;ram[24][68]=0;ram[24][69]=0;ram[24][70]=1;ram[24][71]=0;ram[24][72]=1;ram[24][73]=0;ram[24][74]=1;ram[24][75]=0;ram[24][76]=1;ram[24][77]=0;ram[24][78]=1;ram[24][79]=0;ram[24][80]=1;ram[24][81]=0;ram[24][82]=0;ram[24][83]=0;ram[24][84]=1;ram[24][85]=0;ram[24][86]=1;ram[24][87]=0;ram[24][88]=1;ram[24][89]=0;ram[24][90]=1;ram[24][91]=0;ram[24][92]=0;ram[24][93]=0;ram[24][94]=1;ram[24][95]=0;ram[24][96]=0;ram[24][97]=0;ram[24][98]=0;ram[24][99]=0;ram[24][100]=0;ram[24][101]=0;ram[24][102]=0;ram[24][103]=0;ram[24][104]=0;ram[24][105]=0;ram[24][106]=0;ram[24][107]=0;ram[24][108]=0;ram[24][109]=0;ram[24][110]=0;ram[24][111]=0;ram[24][112]=0;ram[24][113]=0;ram[24][114]=0;ram[24][115]=0;ram[24][116]=0;ram[24][117]=0;ram[24][118]=0;ram[24][119]=0;ram[24][120]=0;ram[24][121]=0;ram[24][122]=0;ram[24][123]=0;ram[24][124]=0;ram[24][125]=0;ram[24][126]=0;ram[24][127]=0;ram[24][128]=0;ram[24][129]=0;ram[24][130]=0;ram[24][131]=0;ram[24][132]=0;ram[24][133]=0;ram[24][134]=0;ram[24][135]=0;ram[24][136]=0;ram[24][137]=0;ram[24][138]=0;ram[24][139]=0;ram[24][140]=0;
        ram[25][0]=0;ram[25][1]=0;ram[25][2]=0;ram[25][3]=0;ram[25][4]=0;ram[25][5]=0;ram[25][6]=0;ram[25][7]=0;ram[25][8]=0;ram[25][9]=0;ram[25][10]=0;ram[25][11]=0;ram[25][12]=0;ram[25][13]=0;ram[25][14]=0;ram[25][15]=0;ram[25][16]=0;ram[25][17]=0;ram[25][18]=0;ram[25][19]=0;ram[25][20]=0;ram[25][21]=0;ram[25][22]=0;ram[25][23]=0;ram[25][24]=0;ram[25][25]=0;ram[25][26]=0;ram[25][27]=0;ram[25][28]=0;ram[25][29]=0;ram[25][30]=0;ram[25][31]=0;ram[25][32]=0;ram[25][33]=0;ram[25][34]=0;ram[25][35]=0;ram[25][36]=0;ram[25][37]=0;ram[25][38]=0;ram[25][39]=0;ram[25][40]=0;ram[25][41]=0;ram[25][42]=0;ram[25][43]=0;ram[25][44]=0;ram[25][45]=1;ram[25][46]=0;ram[25][47]=1;ram[25][48]=0;ram[25][49]=1;ram[25][50]=0;ram[25][51]=1;ram[25][52]=0;ram[25][53]=1;ram[25][54]=0;ram[25][55]=1;ram[25][56]=0;ram[25][57]=0;ram[25][58]=0;ram[25][59]=1;ram[25][60]=0;ram[25][61]=1;ram[25][62]=0;ram[25][63]=1;ram[25][64]=0;ram[25][65]=0;ram[25][66]=0;ram[25][67]=0;ram[25][68]=0;ram[25][69]=1;ram[25][70]=0;ram[25][71]=0;ram[25][72]=0;ram[25][73]=1;ram[25][74]=0;ram[25][75]=1;ram[25][76]=0;ram[25][77]=1;ram[25][78]=0;ram[25][79]=0;ram[25][80]=0;ram[25][81]=1;ram[25][82]=0;ram[25][83]=1;ram[25][84]=0;ram[25][85]=1;ram[25][86]=0;ram[25][87]=0;ram[25][88]=0;ram[25][89]=1;ram[25][90]=0;ram[25][91]=0;ram[25][92]=0;ram[25][93]=1;ram[25][94]=0;ram[25][95]=1;ram[25][96]=0;ram[25][97]=0;ram[25][98]=0;ram[25][99]=0;ram[25][100]=0;ram[25][101]=0;ram[25][102]=0;ram[25][103]=0;ram[25][104]=0;ram[25][105]=0;ram[25][106]=0;ram[25][107]=0;ram[25][108]=0;ram[25][109]=0;ram[25][110]=0;ram[25][111]=0;ram[25][112]=0;ram[25][113]=0;ram[25][114]=0;ram[25][115]=0;ram[25][116]=0;ram[25][117]=0;ram[25][118]=0;ram[25][119]=0;ram[25][120]=0;ram[25][121]=0;ram[25][122]=0;ram[25][123]=0;ram[25][124]=0;ram[25][125]=0;ram[25][126]=0;ram[25][127]=0;ram[25][128]=0;ram[25][129]=0;ram[25][130]=0;ram[25][131]=0;ram[25][132]=0;ram[25][133]=0;ram[25][134]=0;ram[25][135]=0;ram[25][136]=0;ram[25][137]=0;ram[25][138]=0;ram[25][139]=0;ram[25][140]=0;
        ram[26][0]=0;ram[26][1]=0;ram[26][2]=0;ram[26][3]=0;ram[26][4]=0;ram[26][5]=0;ram[26][6]=0;ram[26][7]=0;ram[26][8]=0;ram[26][9]=0;ram[26][10]=0;ram[26][11]=0;ram[26][12]=0;ram[26][13]=0;ram[26][14]=0;ram[26][15]=0;ram[26][16]=0;ram[26][17]=0;ram[26][18]=0;ram[26][19]=0;ram[26][20]=0;ram[26][21]=0;ram[26][22]=0;ram[26][23]=0;ram[26][24]=0;ram[26][25]=0;ram[26][26]=0;ram[26][27]=0;ram[26][28]=0;ram[26][29]=0;ram[26][30]=0;ram[26][31]=0;ram[26][32]=0;ram[26][33]=0;ram[26][34]=0;ram[26][35]=0;ram[26][36]=0;ram[26][37]=0;ram[26][38]=0;ram[26][39]=0;ram[26][40]=0;ram[26][41]=0;ram[26][42]=0;ram[26][43]=0;ram[26][44]=1;ram[26][45]=0;ram[26][46]=0;ram[26][47]=0;ram[26][48]=1;ram[26][49]=0;ram[26][50]=1;ram[26][51]=0;ram[26][52]=1;ram[26][53]=0;ram[26][54]=1;ram[26][55]=0;ram[26][56]=0;ram[26][57]=0;ram[26][58]=1;ram[26][59]=0;ram[26][60]=0;ram[26][61]=0;ram[26][62]=1;ram[26][63]=0;ram[26][64]=0;ram[26][65]=0;ram[26][66]=1;ram[26][67]=0;ram[26][68]=1;ram[26][69]=0;ram[26][70]=1;ram[26][71]=0;ram[26][72]=0;ram[26][73]=0;ram[26][74]=0;ram[26][75]=0;ram[26][76]=1;ram[26][77]=0;ram[26][78]=1;ram[26][79]=0;ram[26][80]=0;ram[26][81]=0;ram[26][82]=0;ram[26][83]=0;ram[26][84]=0;ram[26][85]=0;ram[26][86]=0;ram[26][87]=0;ram[26][88]=1;ram[26][89]=0;ram[26][90]=1;ram[26][91]=0;ram[26][92]=0;ram[26][93]=0;ram[26][94]=0;ram[26][95]=0;ram[26][96]=1;ram[26][97]=0;ram[26][98]=0;ram[26][99]=0;ram[26][100]=0;ram[26][101]=0;ram[26][102]=0;ram[26][103]=0;ram[26][104]=0;ram[26][105]=0;ram[26][106]=0;ram[26][107]=0;ram[26][108]=0;ram[26][109]=0;ram[26][110]=0;ram[26][111]=0;ram[26][112]=0;ram[26][113]=0;ram[26][114]=0;ram[26][115]=0;ram[26][116]=0;ram[26][117]=0;ram[26][118]=0;ram[26][119]=0;ram[26][120]=0;ram[26][121]=0;ram[26][122]=0;ram[26][123]=0;ram[26][124]=0;ram[26][125]=0;ram[26][126]=0;ram[26][127]=0;ram[26][128]=0;ram[26][129]=0;ram[26][130]=0;ram[26][131]=0;ram[26][132]=0;ram[26][133]=0;ram[26][134]=0;ram[26][135]=0;ram[26][136]=0;ram[26][137]=0;ram[26][138]=0;ram[26][139]=0;ram[26][140]=0;
        ram[27][0]=0;ram[27][1]=0;ram[27][2]=0;ram[27][3]=0;ram[27][4]=0;ram[27][5]=0;ram[27][6]=0;ram[27][7]=0;ram[27][8]=0;ram[27][9]=0;ram[27][10]=0;ram[27][11]=0;ram[27][12]=0;ram[27][13]=0;ram[27][14]=0;ram[27][15]=0;ram[27][16]=0;ram[27][17]=0;ram[27][18]=0;ram[27][19]=0;ram[27][20]=0;ram[27][21]=0;ram[27][22]=0;ram[27][23]=0;ram[27][24]=0;ram[27][25]=0;ram[27][26]=0;ram[27][27]=0;ram[27][28]=0;ram[27][29]=0;ram[27][30]=0;ram[27][31]=0;ram[27][32]=0;ram[27][33]=0;ram[27][34]=0;ram[27][35]=0;ram[27][36]=0;ram[27][37]=0;ram[27][38]=0;ram[27][39]=0;ram[27][40]=0;ram[27][41]=0;ram[27][42]=0;ram[27][43]=1;ram[27][44]=0;ram[27][45]=0;ram[27][46]=0;ram[27][47]=1;ram[27][48]=0;ram[27][49]=1;ram[27][50]=0;ram[27][51]=1;ram[27][52]=0;ram[27][53]=1;ram[27][54]=0;ram[27][55]=1;ram[27][56]=0;ram[27][57]=1;ram[27][58]=0;ram[27][59]=1;ram[27][60]=0;ram[27][61]=1;ram[27][62]=0;ram[27][63]=0;ram[27][64]=0;ram[27][65]=1;ram[27][66]=0;ram[27][67]=0;ram[27][68]=0;ram[27][69]=1;ram[27][70]=0;ram[27][71]=1;ram[27][72]=0;ram[27][73]=1;ram[27][74]=0;ram[27][75]=1;ram[27][76]=0;ram[27][77]=0;ram[27][78]=0;ram[27][79]=0;ram[27][80]=0;ram[27][81]=1;ram[27][82]=0;ram[27][83]=1;ram[27][84]=0;ram[27][85]=1;ram[27][86]=0;ram[27][87]=1;ram[27][88]=0;ram[27][89]=1;ram[27][90]=0;ram[27][91]=0;ram[27][92]=0;ram[27][93]=1;ram[27][94]=0;ram[27][95]=0;ram[27][96]=0;ram[27][97]=1;ram[27][98]=0;ram[27][99]=0;ram[27][100]=0;ram[27][101]=0;ram[27][102]=0;ram[27][103]=0;ram[27][104]=0;ram[27][105]=0;ram[27][106]=0;ram[27][107]=0;ram[27][108]=0;ram[27][109]=0;ram[27][110]=0;ram[27][111]=0;ram[27][112]=0;ram[27][113]=0;ram[27][114]=0;ram[27][115]=0;ram[27][116]=0;ram[27][117]=0;ram[27][118]=0;ram[27][119]=0;ram[27][120]=0;ram[27][121]=0;ram[27][122]=0;ram[27][123]=0;ram[27][124]=0;ram[27][125]=0;ram[27][126]=0;ram[27][127]=0;ram[27][128]=0;ram[27][129]=0;ram[27][130]=0;ram[27][131]=0;ram[27][132]=0;ram[27][133]=0;ram[27][134]=0;ram[27][135]=0;ram[27][136]=0;ram[27][137]=0;ram[27][138]=0;ram[27][139]=0;ram[27][140]=0;
        ram[28][0]=0;ram[28][1]=0;ram[28][2]=0;ram[28][3]=0;ram[28][4]=0;ram[28][5]=0;ram[28][6]=0;ram[28][7]=0;ram[28][8]=0;ram[28][9]=0;ram[28][10]=0;ram[28][11]=0;ram[28][12]=0;ram[28][13]=0;ram[28][14]=0;ram[28][15]=0;ram[28][16]=0;ram[28][17]=0;ram[28][18]=0;ram[28][19]=0;ram[28][20]=0;ram[28][21]=0;ram[28][22]=0;ram[28][23]=0;ram[28][24]=0;ram[28][25]=0;ram[28][26]=0;ram[28][27]=0;ram[28][28]=0;ram[28][29]=0;ram[28][30]=0;ram[28][31]=0;ram[28][32]=0;ram[28][33]=0;ram[28][34]=0;ram[28][35]=0;ram[28][36]=0;ram[28][37]=0;ram[28][38]=0;ram[28][39]=0;ram[28][40]=0;ram[28][41]=0;ram[28][42]=1;ram[28][43]=0;ram[28][44]=0;ram[28][45]=0;ram[28][46]=1;ram[28][47]=0;ram[28][48]=1;ram[28][49]=0;ram[28][50]=0;ram[28][51]=0;ram[28][52]=1;ram[28][53]=0;ram[28][54]=0;ram[28][55]=0;ram[28][56]=1;ram[28][57]=0;ram[28][58]=0;ram[28][59]=0;ram[28][60]=1;ram[28][61]=0;ram[28][62]=0;ram[28][63]=0;ram[28][64]=1;ram[28][65]=0;ram[28][66]=1;ram[28][67]=0;ram[28][68]=0;ram[28][69]=0;ram[28][70]=1;ram[28][71]=0;ram[28][72]=0;ram[28][73]=0;ram[28][74]=0;ram[28][75]=0;ram[28][76]=1;ram[28][77]=0;ram[28][78]=1;ram[28][79]=0;ram[28][80]=1;ram[28][81]=0;ram[28][82]=1;ram[28][83]=0;ram[28][84]=0;ram[28][85]=0;ram[28][86]=1;ram[28][87]=0;ram[28][88]=1;ram[28][89]=0;ram[28][90]=1;ram[28][91]=0;ram[28][92]=1;ram[28][93]=0;ram[28][94]=1;ram[28][95]=0;ram[28][96]=1;ram[28][97]=0;ram[28][98]=1;ram[28][99]=0;ram[28][100]=0;ram[28][101]=0;ram[28][102]=0;ram[28][103]=0;ram[28][104]=0;ram[28][105]=0;ram[28][106]=0;ram[28][107]=0;ram[28][108]=0;ram[28][109]=0;ram[28][110]=0;ram[28][111]=0;ram[28][112]=0;ram[28][113]=0;ram[28][114]=0;ram[28][115]=0;ram[28][116]=0;ram[28][117]=0;ram[28][118]=0;ram[28][119]=0;ram[28][120]=0;ram[28][121]=0;ram[28][122]=0;ram[28][123]=0;ram[28][124]=0;ram[28][125]=0;ram[28][126]=0;ram[28][127]=0;ram[28][128]=0;ram[28][129]=0;ram[28][130]=0;ram[28][131]=0;ram[28][132]=0;ram[28][133]=0;ram[28][134]=0;ram[28][135]=0;ram[28][136]=0;ram[28][137]=0;ram[28][138]=0;ram[28][139]=0;ram[28][140]=0;
        ram[29][0]=0;ram[29][1]=0;ram[29][2]=0;ram[29][3]=0;ram[29][4]=0;ram[29][5]=0;ram[29][6]=0;ram[29][7]=0;ram[29][8]=0;ram[29][9]=0;ram[29][10]=0;ram[29][11]=0;ram[29][12]=0;ram[29][13]=0;ram[29][14]=0;ram[29][15]=0;ram[29][16]=0;ram[29][17]=0;ram[29][18]=0;ram[29][19]=0;ram[29][20]=0;ram[29][21]=0;ram[29][22]=0;ram[29][23]=0;ram[29][24]=0;ram[29][25]=0;ram[29][26]=0;ram[29][27]=0;ram[29][28]=0;ram[29][29]=0;ram[29][30]=0;ram[29][31]=0;ram[29][32]=0;ram[29][33]=0;ram[29][34]=0;ram[29][35]=0;ram[29][36]=0;ram[29][37]=0;ram[29][38]=0;ram[29][39]=0;ram[29][40]=0;ram[29][41]=1;ram[29][42]=0;ram[29][43]=0;ram[29][44]=0;ram[29][45]=0;ram[29][46]=0;ram[29][47]=0;ram[29][48]=0;ram[29][49]=0;ram[29][50]=0;ram[29][51]=1;ram[29][52]=0;ram[29][53]=0;ram[29][54]=0;ram[29][55]=1;ram[29][56]=0;ram[29][57]=0;ram[29][58]=0;ram[29][59]=1;ram[29][60]=0;ram[29][61]=0;ram[29][62]=0;ram[29][63]=1;ram[29][64]=0;ram[29][65]=0;ram[29][66]=0;ram[29][67]=1;ram[29][68]=0;ram[29][69]=0;ram[29][70]=0;ram[29][71]=1;ram[29][72]=0;ram[29][73]=1;ram[29][74]=0;ram[29][75]=0;ram[29][76]=0;ram[29][77]=1;ram[29][78]=0;ram[29][79]=1;ram[29][80]=0;ram[29][81]=1;ram[29][82]=0;ram[29][83]=0;ram[29][84]=0;ram[29][85]=0;ram[29][86]=0;ram[29][87]=0;ram[29][88]=0;ram[29][89]=1;ram[29][90]=0;ram[29][91]=0;ram[29][92]=0;ram[29][93]=1;ram[29][94]=0;ram[29][95]=0;ram[29][96]=0;ram[29][97]=1;ram[29][98]=0;ram[29][99]=1;ram[29][100]=0;ram[29][101]=0;ram[29][102]=0;ram[29][103]=0;ram[29][104]=0;ram[29][105]=0;ram[29][106]=0;ram[29][107]=0;ram[29][108]=0;ram[29][109]=0;ram[29][110]=0;ram[29][111]=0;ram[29][112]=0;ram[29][113]=0;ram[29][114]=0;ram[29][115]=0;ram[29][116]=0;ram[29][117]=0;ram[29][118]=0;ram[29][119]=0;ram[29][120]=0;ram[29][121]=0;ram[29][122]=0;ram[29][123]=0;ram[29][124]=0;ram[29][125]=0;ram[29][126]=0;ram[29][127]=0;ram[29][128]=0;ram[29][129]=0;ram[29][130]=0;ram[29][131]=0;ram[29][132]=0;ram[29][133]=0;ram[29][134]=0;ram[29][135]=0;ram[29][136]=0;ram[29][137]=0;ram[29][138]=0;ram[29][139]=0;ram[29][140]=0;
        ram[30][0]=0;ram[30][1]=0;ram[30][2]=0;ram[30][3]=0;ram[30][4]=0;ram[30][5]=0;ram[30][6]=0;ram[30][7]=0;ram[30][8]=0;ram[30][9]=0;ram[30][10]=0;ram[30][11]=0;ram[30][12]=0;ram[30][13]=0;ram[30][14]=0;ram[30][15]=0;ram[30][16]=0;ram[30][17]=0;ram[30][18]=0;ram[30][19]=0;ram[30][20]=0;ram[30][21]=0;ram[30][22]=0;ram[30][23]=0;ram[30][24]=0;ram[30][25]=0;ram[30][26]=0;ram[30][27]=0;ram[30][28]=0;ram[30][29]=0;ram[30][30]=0;ram[30][31]=0;ram[30][32]=0;ram[30][33]=0;ram[30][34]=0;ram[30][35]=0;ram[30][36]=0;ram[30][37]=0;ram[30][38]=0;ram[30][39]=0;ram[30][40]=1;ram[30][41]=0;ram[30][42]=1;ram[30][43]=0;ram[30][44]=1;ram[30][45]=0;ram[30][46]=1;ram[30][47]=0;ram[30][48]=1;ram[30][49]=0;ram[30][50]=0;ram[30][51]=0;ram[30][52]=1;ram[30][53]=0;ram[30][54]=0;ram[30][55]=0;ram[30][56]=1;ram[30][57]=0;ram[30][58]=1;ram[30][59]=0;ram[30][60]=1;ram[30][61]=0;ram[30][62]=0;ram[30][63]=0;ram[30][64]=0;ram[30][65]=0;ram[30][66]=1;ram[30][67]=0;ram[30][68]=0;ram[30][69]=0;ram[30][70]=1;ram[30][71]=0;ram[30][72]=1;ram[30][73]=0;ram[30][74]=0;ram[30][75]=0;ram[30][76]=1;ram[30][77]=0;ram[30][78]=0;ram[30][79]=0;ram[30][80]=1;ram[30][81]=0;ram[30][82]=0;ram[30][83]=0;ram[30][84]=1;ram[30][85]=0;ram[30][86]=0;ram[30][87]=0;ram[30][88]=0;ram[30][89]=0;ram[30][90]=1;ram[30][91]=0;ram[30][92]=1;ram[30][93]=0;ram[30][94]=0;ram[30][95]=0;ram[30][96]=1;ram[30][97]=0;ram[30][98]=1;ram[30][99]=0;ram[30][100]=1;ram[30][101]=0;ram[30][102]=0;ram[30][103]=0;ram[30][104]=0;ram[30][105]=0;ram[30][106]=0;ram[30][107]=0;ram[30][108]=0;ram[30][109]=0;ram[30][110]=0;ram[30][111]=0;ram[30][112]=0;ram[30][113]=0;ram[30][114]=0;ram[30][115]=0;ram[30][116]=0;ram[30][117]=0;ram[30][118]=0;ram[30][119]=0;ram[30][120]=0;ram[30][121]=0;ram[30][122]=0;ram[30][123]=0;ram[30][124]=0;ram[30][125]=0;ram[30][126]=0;ram[30][127]=0;ram[30][128]=0;ram[30][129]=0;ram[30][130]=0;ram[30][131]=0;ram[30][132]=0;ram[30][133]=0;ram[30][134]=0;ram[30][135]=0;ram[30][136]=0;ram[30][137]=0;ram[30][138]=0;ram[30][139]=0;ram[30][140]=0;
        ram[31][0]=0;ram[31][1]=0;ram[31][2]=0;ram[31][3]=0;ram[31][4]=0;ram[31][5]=0;ram[31][6]=0;ram[31][7]=0;ram[31][8]=0;ram[31][9]=0;ram[31][10]=0;ram[31][11]=0;ram[31][12]=0;ram[31][13]=0;ram[31][14]=0;ram[31][15]=0;ram[31][16]=0;ram[31][17]=0;ram[31][18]=0;ram[31][19]=0;ram[31][20]=0;ram[31][21]=0;ram[31][22]=0;ram[31][23]=0;ram[31][24]=0;ram[31][25]=0;ram[31][26]=0;ram[31][27]=0;ram[31][28]=0;ram[31][29]=0;ram[31][30]=0;ram[31][31]=0;ram[31][32]=0;ram[31][33]=0;ram[31][34]=0;ram[31][35]=0;ram[31][36]=0;ram[31][37]=0;ram[31][38]=0;ram[31][39]=1;ram[31][40]=0;ram[31][41]=0;ram[31][42]=0;ram[31][43]=0;ram[31][44]=0;ram[31][45]=1;ram[31][46]=0;ram[31][47]=1;ram[31][48]=0;ram[31][49]=1;ram[31][50]=0;ram[31][51]=0;ram[31][52]=0;ram[31][53]=1;ram[31][54]=0;ram[31][55]=1;ram[31][56]=0;ram[31][57]=0;ram[31][58]=0;ram[31][59]=0;ram[31][60]=0;ram[31][61]=0;ram[31][62]=0;ram[31][63]=1;ram[31][64]=0;ram[31][65]=1;ram[31][66]=0;ram[31][67]=0;ram[31][68]=0;ram[31][69]=1;ram[31][70]=0;ram[31][71]=0;ram[31][72]=0;ram[31][73]=1;ram[31][74]=0;ram[31][75]=1;ram[31][76]=0;ram[31][77]=1;ram[31][78]=0;ram[31][79]=1;ram[31][80]=0;ram[31][81]=0;ram[31][82]=0;ram[31][83]=0;ram[31][84]=0;ram[31][85]=0;ram[31][86]=0;ram[31][87]=1;ram[31][88]=0;ram[31][89]=0;ram[31][90]=0;ram[31][91]=1;ram[31][92]=0;ram[31][93]=1;ram[31][94]=0;ram[31][95]=1;ram[31][96]=0;ram[31][97]=1;ram[31][98]=0;ram[31][99]=1;ram[31][100]=0;ram[31][101]=1;ram[31][102]=0;ram[31][103]=0;ram[31][104]=0;ram[31][105]=0;ram[31][106]=0;ram[31][107]=0;ram[31][108]=0;ram[31][109]=0;ram[31][110]=0;ram[31][111]=0;ram[31][112]=0;ram[31][113]=0;ram[31][114]=0;ram[31][115]=0;ram[31][116]=0;ram[31][117]=0;ram[31][118]=0;ram[31][119]=0;ram[31][120]=0;ram[31][121]=0;ram[31][122]=0;ram[31][123]=0;ram[31][124]=0;ram[31][125]=0;ram[31][126]=0;ram[31][127]=0;ram[31][128]=0;ram[31][129]=0;ram[31][130]=0;ram[31][131]=0;ram[31][132]=0;ram[31][133]=0;ram[31][134]=0;ram[31][135]=0;ram[31][136]=0;ram[31][137]=0;ram[31][138]=0;ram[31][139]=0;ram[31][140]=0;
        ram[32][0]=0;ram[32][1]=0;ram[32][2]=0;ram[32][3]=0;ram[32][4]=0;ram[32][5]=0;ram[32][6]=0;ram[32][7]=0;ram[32][8]=0;ram[32][9]=0;ram[32][10]=0;ram[32][11]=0;ram[32][12]=0;ram[32][13]=0;ram[32][14]=0;ram[32][15]=0;ram[32][16]=0;ram[32][17]=0;ram[32][18]=0;ram[32][19]=0;ram[32][20]=0;ram[32][21]=0;ram[32][22]=0;ram[32][23]=0;ram[32][24]=0;ram[32][25]=0;ram[32][26]=0;ram[32][27]=0;ram[32][28]=0;ram[32][29]=0;ram[32][30]=0;ram[32][31]=0;ram[32][32]=0;ram[32][33]=0;ram[32][34]=0;ram[32][35]=0;ram[32][36]=0;ram[32][37]=0;ram[32][38]=1;ram[32][39]=0;ram[32][40]=1;ram[32][41]=0;ram[32][42]=1;ram[32][43]=0;ram[32][44]=1;ram[32][45]=0;ram[32][46]=1;ram[32][47]=0;ram[32][48]=0;ram[32][49]=0;ram[32][50]=1;ram[32][51]=0;ram[32][52]=0;ram[32][53]=0;ram[32][54]=1;ram[32][55]=0;ram[32][56]=1;ram[32][57]=0;ram[32][58]=1;ram[32][59]=0;ram[32][60]=1;ram[32][61]=0;ram[32][62]=1;ram[32][63]=0;ram[32][64]=0;ram[32][65]=0;ram[32][66]=1;ram[32][67]=0;ram[32][68]=1;ram[32][69]=0;ram[32][70]=1;ram[32][71]=0;ram[32][72]=0;ram[32][73]=0;ram[32][74]=0;ram[32][75]=0;ram[32][76]=0;ram[32][77]=0;ram[32][78]=1;ram[32][79]=0;ram[32][80]=1;ram[32][81]=0;ram[32][82]=0;ram[32][83]=0;ram[32][84]=0;ram[32][85]=0;ram[32][86]=1;ram[32][87]=0;ram[32][88]=1;ram[32][89]=0;ram[32][90]=1;ram[32][91]=0;ram[32][92]=0;ram[32][93]=0;ram[32][94]=0;ram[32][95]=0;ram[32][96]=1;ram[32][97]=0;ram[32][98]=1;ram[32][99]=0;ram[32][100]=1;ram[32][101]=0;ram[32][102]=1;ram[32][103]=0;ram[32][104]=0;ram[32][105]=0;ram[32][106]=0;ram[32][107]=0;ram[32][108]=0;ram[32][109]=0;ram[32][110]=0;ram[32][111]=0;ram[32][112]=0;ram[32][113]=0;ram[32][114]=0;ram[32][115]=0;ram[32][116]=0;ram[32][117]=0;ram[32][118]=0;ram[32][119]=0;ram[32][120]=0;ram[32][121]=0;ram[32][122]=0;ram[32][123]=0;ram[32][124]=0;ram[32][125]=0;ram[32][126]=0;ram[32][127]=0;ram[32][128]=0;ram[32][129]=0;ram[32][130]=0;ram[32][131]=0;ram[32][132]=0;ram[32][133]=0;ram[32][134]=0;ram[32][135]=0;ram[32][136]=0;ram[32][137]=0;ram[32][138]=0;ram[32][139]=0;ram[32][140]=0;
        ram[33][0]=0;ram[33][1]=0;ram[33][2]=0;ram[33][3]=0;ram[33][4]=0;ram[33][5]=0;ram[33][6]=0;ram[33][7]=0;ram[33][8]=0;ram[33][9]=0;ram[33][10]=0;ram[33][11]=0;ram[33][12]=0;ram[33][13]=0;ram[33][14]=0;ram[33][15]=0;ram[33][16]=0;ram[33][17]=0;ram[33][18]=0;ram[33][19]=0;ram[33][20]=0;ram[33][21]=0;ram[33][22]=0;ram[33][23]=0;ram[33][24]=0;ram[33][25]=0;ram[33][26]=0;ram[33][27]=0;ram[33][28]=0;ram[33][29]=0;ram[33][30]=0;ram[33][31]=0;ram[33][32]=0;ram[33][33]=0;ram[33][34]=0;ram[33][35]=0;ram[33][36]=0;ram[33][37]=1;ram[33][38]=0;ram[33][39]=1;ram[33][40]=0;ram[33][41]=1;ram[33][42]=0;ram[33][43]=1;ram[33][44]=0;ram[33][45]=1;ram[33][46]=0;ram[33][47]=1;ram[33][48]=0;ram[33][49]=0;ram[33][50]=0;ram[33][51]=0;ram[33][52]=0;ram[33][53]=1;ram[33][54]=0;ram[33][55]=1;ram[33][56]=0;ram[33][57]=1;ram[33][58]=0;ram[33][59]=1;ram[33][60]=0;ram[33][61]=0;ram[33][62]=0;ram[33][63]=0;ram[33][64]=0;ram[33][65]=0;ram[33][66]=0;ram[33][67]=1;ram[33][68]=0;ram[33][69]=0;ram[33][70]=0;ram[33][71]=1;ram[33][72]=0;ram[33][73]=0;ram[33][74]=0;ram[33][75]=1;ram[33][76]=0;ram[33][77]=1;ram[33][78]=0;ram[33][79]=1;ram[33][80]=0;ram[33][81]=0;ram[33][82]=0;ram[33][83]=1;ram[33][84]=0;ram[33][85]=1;ram[33][86]=0;ram[33][87]=1;ram[33][88]=0;ram[33][89]=1;ram[33][90]=0;ram[33][91]=1;ram[33][92]=0;ram[33][93]=1;ram[33][94]=0;ram[33][95]=0;ram[33][96]=0;ram[33][97]=1;ram[33][98]=0;ram[33][99]=1;ram[33][100]=0;ram[33][101]=1;ram[33][102]=0;ram[33][103]=1;ram[33][104]=0;ram[33][105]=0;ram[33][106]=0;ram[33][107]=0;ram[33][108]=0;ram[33][109]=0;ram[33][110]=0;ram[33][111]=0;ram[33][112]=0;ram[33][113]=0;ram[33][114]=0;ram[33][115]=0;ram[33][116]=0;ram[33][117]=0;ram[33][118]=0;ram[33][119]=0;ram[33][120]=0;ram[33][121]=0;ram[33][122]=0;ram[33][123]=0;ram[33][124]=0;ram[33][125]=0;ram[33][126]=0;ram[33][127]=0;ram[33][128]=0;ram[33][129]=0;ram[33][130]=0;ram[33][131]=0;ram[33][132]=0;ram[33][133]=0;ram[33][134]=0;ram[33][135]=0;ram[33][136]=0;ram[33][137]=0;ram[33][138]=0;ram[33][139]=0;ram[33][140]=0;
        ram[34][0]=0;ram[34][1]=0;ram[34][2]=0;ram[34][3]=0;ram[34][4]=0;ram[34][5]=0;ram[34][6]=0;ram[34][7]=0;ram[34][8]=0;ram[34][9]=0;ram[34][10]=0;ram[34][11]=0;ram[34][12]=0;ram[34][13]=0;ram[34][14]=0;ram[34][15]=0;ram[34][16]=0;ram[34][17]=0;ram[34][18]=0;ram[34][19]=0;ram[34][20]=0;ram[34][21]=0;ram[34][22]=0;ram[34][23]=0;ram[34][24]=0;ram[34][25]=0;ram[34][26]=0;ram[34][27]=0;ram[34][28]=0;ram[34][29]=0;ram[34][30]=0;ram[34][31]=0;ram[34][32]=0;ram[34][33]=0;ram[34][34]=0;ram[34][35]=0;ram[34][36]=1;ram[34][37]=0;ram[34][38]=0;ram[34][39]=0;ram[34][40]=1;ram[34][41]=0;ram[34][42]=1;ram[34][43]=0;ram[34][44]=1;ram[34][45]=0;ram[34][46]=1;ram[34][47]=0;ram[34][48]=1;ram[34][49]=0;ram[34][50]=0;ram[34][51]=0;ram[34][52]=0;ram[34][53]=0;ram[34][54]=1;ram[34][55]=0;ram[34][56]=0;ram[34][57]=0;ram[34][58]=1;ram[34][59]=0;ram[34][60]=0;ram[34][61]=0;ram[34][62]=0;ram[34][63]=0;ram[34][64]=1;ram[34][65]=0;ram[34][66]=1;ram[34][67]=0;ram[34][68]=0;ram[34][69]=0;ram[34][70]=0;ram[34][71]=0;ram[34][72]=1;ram[34][73]=0;ram[34][74]=1;ram[34][75]=0;ram[34][76]=1;ram[34][77]=0;ram[34][78]=1;ram[34][79]=0;ram[34][80]=1;ram[34][81]=0;ram[34][82]=1;ram[34][83]=0;ram[34][84]=1;ram[34][85]=0;ram[34][86]=1;ram[34][87]=0;ram[34][88]=0;ram[34][89]=0;ram[34][90]=1;ram[34][91]=0;ram[34][92]=0;ram[34][93]=0;ram[34][94]=0;ram[34][95]=0;ram[34][96]=1;ram[34][97]=0;ram[34][98]=1;ram[34][99]=0;ram[34][100]=1;ram[34][101]=0;ram[34][102]=1;ram[34][103]=0;ram[34][104]=1;ram[34][105]=0;ram[34][106]=0;ram[34][107]=0;ram[34][108]=0;ram[34][109]=0;ram[34][110]=0;ram[34][111]=0;ram[34][112]=0;ram[34][113]=0;ram[34][114]=0;ram[34][115]=0;ram[34][116]=0;ram[34][117]=0;ram[34][118]=0;ram[34][119]=0;ram[34][120]=0;ram[34][121]=0;ram[34][122]=0;ram[34][123]=0;ram[34][124]=0;ram[34][125]=0;ram[34][126]=0;ram[34][127]=0;ram[34][128]=0;ram[34][129]=0;ram[34][130]=0;ram[34][131]=0;ram[34][132]=0;ram[34][133]=0;ram[34][134]=0;ram[34][135]=0;ram[34][136]=0;ram[34][137]=0;ram[34][138]=0;ram[34][139]=0;ram[34][140]=0;
        ram[35][0]=0;ram[35][1]=0;ram[35][2]=0;ram[35][3]=0;ram[35][4]=0;ram[35][5]=0;ram[35][6]=0;ram[35][7]=0;ram[35][8]=0;ram[35][9]=0;ram[35][10]=0;ram[35][11]=0;ram[35][12]=0;ram[35][13]=0;ram[35][14]=0;ram[35][15]=0;ram[35][16]=0;ram[35][17]=0;ram[35][18]=0;ram[35][19]=0;ram[35][20]=0;ram[35][21]=0;ram[35][22]=0;ram[35][23]=0;ram[35][24]=0;ram[35][25]=0;ram[35][26]=0;ram[35][27]=0;ram[35][28]=0;ram[35][29]=0;ram[35][30]=0;ram[35][31]=0;ram[35][32]=0;ram[35][33]=0;ram[35][34]=0;ram[35][35]=1;ram[35][36]=0;ram[35][37]=0;ram[35][38]=0;ram[35][39]=1;ram[35][40]=0;ram[35][41]=0;ram[35][42]=0;ram[35][43]=1;ram[35][44]=0;ram[35][45]=0;ram[35][46]=0;ram[35][47]=1;ram[35][48]=0;ram[35][49]=1;ram[35][50]=0;ram[35][51]=0;ram[35][52]=0;ram[35][53]=1;ram[35][54]=0;ram[35][55]=1;ram[35][56]=0;ram[35][57]=1;ram[35][58]=0;ram[35][59]=1;ram[35][60]=0;ram[35][61]=0;ram[35][62]=0;ram[35][63]=1;ram[35][64]=0;ram[35][65]=0;ram[35][66]=0;ram[35][67]=1;ram[35][68]=0;ram[35][69]=0;ram[35][70]=0;ram[35][71]=0;ram[35][72]=0;ram[35][73]=0;ram[35][74]=0;ram[35][75]=1;ram[35][76]=0;ram[35][77]=1;ram[35][78]=0;ram[35][79]=0;ram[35][80]=0;ram[35][81]=1;ram[35][82]=0;ram[35][83]=1;ram[35][84]=0;ram[35][85]=1;ram[35][86]=0;ram[35][87]=1;ram[35][88]=0;ram[35][89]=1;ram[35][90]=0;ram[35][91]=0;ram[35][92]=0;ram[35][93]=1;ram[35][94]=0;ram[35][95]=1;ram[35][96]=0;ram[35][97]=0;ram[35][98]=0;ram[35][99]=0;ram[35][100]=0;ram[35][101]=1;ram[35][102]=0;ram[35][103]=0;ram[35][104]=0;ram[35][105]=1;ram[35][106]=0;ram[35][107]=0;ram[35][108]=0;ram[35][109]=0;ram[35][110]=0;ram[35][111]=0;ram[35][112]=0;ram[35][113]=0;ram[35][114]=0;ram[35][115]=0;ram[35][116]=0;ram[35][117]=0;ram[35][118]=0;ram[35][119]=0;ram[35][120]=0;ram[35][121]=0;ram[35][122]=0;ram[35][123]=0;ram[35][124]=0;ram[35][125]=0;ram[35][126]=0;ram[35][127]=0;ram[35][128]=0;ram[35][129]=0;ram[35][130]=0;ram[35][131]=0;ram[35][132]=0;ram[35][133]=0;ram[35][134]=0;ram[35][135]=0;ram[35][136]=0;ram[35][137]=0;ram[35][138]=0;ram[35][139]=0;ram[35][140]=0;
        ram[36][0]=0;ram[36][1]=0;ram[36][2]=0;ram[36][3]=0;ram[36][4]=0;ram[36][5]=0;ram[36][6]=0;ram[36][7]=0;ram[36][8]=0;ram[36][9]=0;ram[36][10]=0;ram[36][11]=0;ram[36][12]=0;ram[36][13]=0;ram[36][14]=0;ram[36][15]=0;ram[36][16]=0;ram[36][17]=0;ram[36][18]=0;ram[36][19]=0;ram[36][20]=0;ram[36][21]=0;ram[36][22]=0;ram[36][23]=0;ram[36][24]=0;ram[36][25]=0;ram[36][26]=0;ram[36][27]=0;ram[36][28]=0;ram[36][29]=0;ram[36][30]=0;ram[36][31]=0;ram[36][32]=0;ram[36][33]=0;ram[36][34]=1;ram[36][35]=0;ram[36][36]=1;ram[36][37]=0;ram[36][38]=1;ram[36][39]=0;ram[36][40]=1;ram[36][41]=0;ram[36][42]=1;ram[36][43]=0;ram[36][44]=1;ram[36][45]=0;ram[36][46]=0;ram[36][47]=0;ram[36][48]=0;ram[36][49]=0;ram[36][50]=1;ram[36][51]=0;ram[36][52]=1;ram[36][53]=0;ram[36][54]=1;ram[36][55]=0;ram[36][56]=1;ram[36][57]=0;ram[36][58]=1;ram[36][59]=0;ram[36][60]=0;ram[36][61]=0;ram[36][62]=1;ram[36][63]=0;ram[36][64]=0;ram[36][65]=0;ram[36][66]=1;ram[36][67]=0;ram[36][68]=0;ram[36][69]=0;ram[36][70]=0;ram[36][71]=0;ram[36][72]=0;ram[36][73]=0;ram[36][74]=1;ram[36][75]=0;ram[36][76]=1;ram[36][77]=0;ram[36][78]=0;ram[36][79]=0;ram[36][80]=1;ram[36][81]=0;ram[36][82]=0;ram[36][83]=0;ram[36][84]=1;ram[36][85]=0;ram[36][86]=1;ram[36][87]=0;ram[36][88]=1;ram[36][89]=0;ram[36][90]=1;ram[36][91]=0;ram[36][92]=1;ram[36][93]=0;ram[36][94]=1;ram[36][95]=0;ram[36][96]=1;ram[36][97]=0;ram[36][98]=1;ram[36][99]=0;ram[36][100]=0;ram[36][101]=0;ram[36][102]=1;ram[36][103]=0;ram[36][104]=1;ram[36][105]=0;ram[36][106]=1;ram[36][107]=0;ram[36][108]=0;ram[36][109]=0;ram[36][110]=0;ram[36][111]=0;ram[36][112]=0;ram[36][113]=0;ram[36][114]=0;ram[36][115]=0;ram[36][116]=0;ram[36][117]=0;ram[36][118]=0;ram[36][119]=0;ram[36][120]=0;ram[36][121]=0;ram[36][122]=0;ram[36][123]=0;ram[36][124]=0;ram[36][125]=0;ram[36][126]=0;ram[36][127]=0;ram[36][128]=0;ram[36][129]=0;ram[36][130]=0;ram[36][131]=0;ram[36][132]=0;ram[36][133]=0;ram[36][134]=0;ram[36][135]=0;ram[36][136]=0;ram[36][137]=0;ram[36][138]=0;ram[36][139]=0;ram[36][140]=0;
        ram[37][0]=0;ram[37][1]=0;ram[37][2]=0;ram[37][3]=0;ram[37][4]=0;ram[37][5]=0;ram[37][6]=0;ram[37][7]=0;ram[37][8]=0;ram[37][9]=0;ram[37][10]=0;ram[37][11]=0;ram[37][12]=0;ram[37][13]=0;ram[37][14]=0;ram[37][15]=0;ram[37][16]=0;ram[37][17]=0;ram[37][18]=0;ram[37][19]=0;ram[37][20]=0;ram[37][21]=0;ram[37][22]=0;ram[37][23]=0;ram[37][24]=0;ram[37][25]=0;ram[37][26]=0;ram[37][27]=0;ram[37][28]=0;ram[37][29]=0;ram[37][30]=0;ram[37][31]=0;ram[37][32]=0;ram[37][33]=1;ram[37][34]=0;ram[37][35]=1;ram[37][36]=0;ram[37][37]=0;ram[37][38]=0;ram[37][39]=1;ram[37][40]=0;ram[37][41]=0;ram[37][42]=0;ram[37][43]=0;ram[37][44]=0;ram[37][45]=0;ram[37][46]=0;ram[37][47]=0;ram[37][48]=0;ram[37][49]=1;ram[37][50]=0;ram[37][51]=0;ram[37][52]=0;ram[37][53]=0;ram[37][54]=0;ram[37][55]=1;ram[37][56]=0;ram[37][57]=1;ram[37][58]=0;ram[37][59]=0;ram[37][60]=0;ram[37][61]=0;ram[37][62]=0;ram[37][63]=1;ram[37][64]=0;ram[37][65]=0;ram[37][66]=0;ram[37][67]=0;ram[37][68]=0;ram[37][69]=1;ram[37][70]=0;ram[37][71]=1;ram[37][72]=0;ram[37][73]=1;ram[37][74]=0;ram[37][75]=1;ram[37][76]=0;ram[37][77]=1;ram[37][78]=0;ram[37][79]=1;ram[37][80]=0;ram[37][81]=0;ram[37][82]=0;ram[37][83]=0;ram[37][84]=0;ram[37][85]=0;ram[37][86]=0;ram[37][87]=1;ram[37][88]=0;ram[37][89]=0;ram[37][90]=0;ram[37][91]=1;ram[37][92]=0;ram[37][93]=1;ram[37][94]=0;ram[37][95]=1;ram[37][96]=0;ram[37][97]=0;ram[37][98]=0;ram[37][99]=1;ram[37][100]=0;ram[37][101]=1;ram[37][102]=0;ram[37][103]=1;ram[37][104]=0;ram[37][105]=0;ram[37][106]=0;ram[37][107]=1;ram[37][108]=0;ram[37][109]=0;ram[37][110]=0;ram[37][111]=0;ram[37][112]=0;ram[37][113]=0;ram[37][114]=0;ram[37][115]=0;ram[37][116]=0;ram[37][117]=0;ram[37][118]=0;ram[37][119]=0;ram[37][120]=0;ram[37][121]=0;ram[37][122]=0;ram[37][123]=0;ram[37][124]=0;ram[37][125]=0;ram[37][126]=0;ram[37][127]=0;ram[37][128]=0;ram[37][129]=0;ram[37][130]=0;ram[37][131]=0;ram[37][132]=0;ram[37][133]=0;ram[37][134]=0;ram[37][135]=0;ram[37][136]=0;ram[37][137]=0;ram[37][138]=0;ram[37][139]=0;ram[37][140]=0;
        ram[38][0]=0;ram[38][1]=0;ram[38][2]=0;ram[38][3]=0;ram[38][4]=0;ram[38][5]=0;ram[38][6]=0;ram[38][7]=0;ram[38][8]=0;ram[38][9]=0;ram[38][10]=0;ram[38][11]=0;ram[38][12]=0;ram[38][13]=0;ram[38][14]=0;ram[38][15]=0;ram[38][16]=0;ram[38][17]=0;ram[38][18]=0;ram[38][19]=0;ram[38][20]=0;ram[38][21]=0;ram[38][22]=0;ram[38][23]=0;ram[38][24]=0;ram[38][25]=0;ram[38][26]=0;ram[38][27]=0;ram[38][28]=0;ram[38][29]=0;ram[38][30]=0;ram[38][31]=0;ram[38][32]=1;ram[38][33]=0;ram[38][34]=1;ram[38][35]=0;ram[38][36]=1;ram[38][37]=0;ram[38][38]=0;ram[38][39]=0;ram[38][40]=0;ram[38][41]=0;ram[38][42]=1;ram[38][43]=0;ram[38][44]=1;ram[38][45]=0;ram[38][46]=0;ram[38][47]=0;ram[38][48]=1;ram[38][49]=0;ram[38][50]=0;ram[38][51]=0;ram[38][52]=1;ram[38][53]=0;ram[38][54]=1;ram[38][55]=0;ram[38][56]=0;ram[38][57]=0;ram[38][58]=0;ram[38][59]=0;ram[38][60]=1;ram[38][61]=0;ram[38][62]=0;ram[38][63]=0;ram[38][64]=1;ram[38][65]=0;ram[38][66]=0;ram[38][67]=0;ram[38][68]=1;ram[38][69]=0;ram[38][70]=0;ram[38][71]=0;ram[38][72]=1;ram[38][73]=0;ram[38][74]=0;ram[38][75]=0;ram[38][76]=0;ram[38][77]=0;ram[38][78]=1;ram[38][79]=0;ram[38][80]=1;ram[38][81]=0;ram[38][82]=1;ram[38][83]=0;ram[38][84]=1;ram[38][85]=0;ram[38][86]=0;ram[38][87]=0;ram[38][88]=1;ram[38][89]=0;ram[38][90]=1;ram[38][91]=0;ram[38][92]=1;ram[38][93]=0;ram[38][94]=0;ram[38][95]=0;ram[38][96]=1;ram[38][97]=0;ram[38][98]=0;ram[38][99]=0;ram[38][100]=1;ram[38][101]=0;ram[38][102]=1;ram[38][103]=0;ram[38][104]=1;ram[38][105]=0;ram[38][106]=1;ram[38][107]=0;ram[38][108]=1;ram[38][109]=0;ram[38][110]=0;ram[38][111]=0;ram[38][112]=0;ram[38][113]=0;ram[38][114]=0;ram[38][115]=0;ram[38][116]=0;ram[38][117]=0;ram[38][118]=0;ram[38][119]=0;ram[38][120]=0;ram[38][121]=0;ram[38][122]=0;ram[38][123]=0;ram[38][124]=0;ram[38][125]=0;ram[38][126]=0;ram[38][127]=0;ram[38][128]=0;ram[38][129]=0;ram[38][130]=0;ram[38][131]=0;ram[38][132]=0;ram[38][133]=0;ram[38][134]=0;ram[38][135]=0;ram[38][136]=0;ram[38][137]=0;ram[38][138]=0;ram[38][139]=0;ram[38][140]=0;
        ram[39][0]=0;ram[39][1]=0;ram[39][2]=0;ram[39][3]=0;ram[39][4]=0;ram[39][5]=0;ram[39][6]=0;ram[39][7]=0;ram[39][8]=0;ram[39][9]=0;ram[39][10]=0;ram[39][11]=0;ram[39][12]=0;ram[39][13]=0;ram[39][14]=0;ram[39][15]=0;ram[39][16]=0;ram[39][17]=0;ram[39][18]=0;ram[39][19]=0;ram[39][20]=0;ram[39][21]=0;ram[39][22]=0;ram[39][23]=0;ram[39][24]=0;ram[39][25]=0;ram[39][26]=0;ram[39][27]=0;ram[39][28]=0;ram[39][29]=0;ram[39][30]=0;ram[39][31]=1;ram[39][32]=0;ram[39][33]=1;ram[39][34]=0;ram[39][35]=1;ram[39][36]=0;ram[39][37]=0;ram[39][38]=0;ram[39][39]=1;ram[39][40]=0;ram[39][41]=1;ram[39][42]=0;ram[39][43]=0;ram[39][44]=0;ram[39][45]=1;ram[39][46]=0;ram[39][47]=0;ram[39][48]=0;ram[39][49]=1;ram[39][50]=0;ram[39][51]=1;ram[39][52]=0;ram[39][53]=1;ram[39][54]=0;ram[39][55]=1;ram[39][56]=0;ram[39][57]=1;ram[39][58]=0;ram[39][59]=1;ram[39][60]=0;ram[39][61]=1;ram[39][62]=0;ram[39][63]=1;ram[39][64]=0;ram[39][65]=1;ram[39][66]=0;ram[39][67]=1;ram[39][68]=0;ram[39][69]=1;ram[39][70]=0;ram[39][71]=0;ram[39][72]=0;ram[39][73]=0;ram[39][74]=0;ram[39][75]=0;ram[39][76]=0;ram[39][77]=0;ram[39][78]=0;ram[39][79]=0;ram[39][80]=0;ram[39][81]=0;ram[39][82]=0;ram[39][83]=1;ram[39][84]=0;ram[39][85]=1;ram[39][86]=0;ram[39][87]=0;ram[39][88]=0;ram[39][89]=0;ram[39][90]=0;ram[39][91]=1;ram[39][92]=0;ram[39][93]=1;ram[39][94]=0;ram[39][95]=0;ram[39][96]=0;ram[39][97]=1;ram[39][98]=0;ram[39][99]=0;ram[39][100]=0;ram[39][101]=1;ram[39][102]=0;ram[39][103]=1;ram[39][104]=0;ram[39][105]=1;ram[39][106]=0;ram[39][107]=1;ram[39][108]=0;ram[39][109]=1;ram[39][110]=0;ram[39][111]=0;ram[39][112]=0;ram[39][113]=0;ram[39][114]=0;ram[39][115]=0;ram[39][116]=0;ram[39][117]=0;ram[39][118]=0;ram[39][119]=0;ram[39][120]=0;ram[39][121]=0;ram[39][122]=0;ram[39][123]=0;ram[39][124]=0;ram[39][125]=0;ram[39][126]=0;ram[39][127]=0;ram[39][128]=0;ram[39][129]=0;ram[39][130]=0;ram[39][131]=0;ram[39][132]=0;ram[39][133]=0;ram[39][134]=0;ram[39][135]=0;ram[39][136]=0;ram[39][137]=0;ram[39][138]=0;ram[39][139]=0;ram[39][140]=0;
        ram[40][0]=0;ram[40][1]=0;ram[40][2]=0;ram[40][3]=0;ram[40][4]=0;ram[40][5]=0;ram[40][6]=0;ram[40][7]=0;ram[40][8]=0;ram[40][9]=0;ram[40][10]=0;ram[40][11]=0;ram[40][12]=0;ram[40][13]=0;ram[40][14]=0;ram[40][15]=0;ram[40][16]=0;ram[40][17]=0;ram[40][18]=0;ram[40][19]=0;ram[40][20]=0;ram[40][21]=0;ram[40][22]=0;ram[40][23]=0;ram[40][24]=0;ram[40][25]=0;ram[40][26]=0;ram[40][27]=0;ram[40][28]=0;ram[40][29]=0;ram[40][30]=1;ram[40][31]=0;ram[40][32]=0;ram[40][33]=0;ram[40][34]=0;ram[40][35]=0;ram[40][36]=0;ram[40][37]=0;ram[40][38]=1;ram[40][39]=0;ram[40][40]=1;ram[40][41]=0;ram[40][42]=1;ram[40][43]=0;ram[40][44]=1;ram[40][45]=0;ram[40][46]=0;ram[40][47]=0;ram[40][48]=1;ram[40][49]=0;ram[40][50]=1;ram[40][51]=0;ram[40][52]=1;ram[40][53]=0;ram[40][54]=1;ram[40][55]=0;ram[40][56]=0;ram[40][57]=0;ram[40][58]=0;ram[40][59]=0;ram[40][60]=1;ram[40][61]=0;ram[40][62]=1;ram[40][63]=0;ram[40][64]=1;ram[40][65]=0;ram[40][66]=1;ram[40][67]=0;ram[40][68]=1;ram[40][69]=0;ram[40][70]=0;ram[40][71]=0;ram[40][72]=1;ram[40][73]=0;ram[40][74]=0;ram[40][75]=0;ram[40][76]=0;ram[40][77]=0;ram[40][78]=1;ram[40][79]=0;ram[40][80]=1;ram[40][81]=0;ram[40][82]=0;ram[40][83]=0;ram[40][84]=1;ram[40][85]=0;ram[40][86]=0;ram[40][87]=0;ram[40][88]=1;ram[40][89]=0;ram[40][90]=1;ram[40][91]=0;ram[40][92]=1;ram[40][93]=0;ram[40][94]=1;ram[40][95]=0;ram[40][96]=1;ram[40][97]=0;ram[40][98]=1;ram[40][99]=0;ram[40][100]=1;ram[40][101]=0;ram[40][102]=0;ram[40][103]=0;ram[40][104]=0;ram[40][105]=0;ram[40][106]=1;ram[40][107]=0;ram[40][108]=1;ram[40][109]=0;ram[40][110]=1;ram[40][111]=0;ram[40][112]=0;ram[40][113]=0;ram[40][114]=0;ram[40][115]=0;ram[40][116]=0;ram[40][117]=0;ram[40][118]=0;ram[40][119]=0;ram[40][120]=0;ram[40][121]=0;ram[40][122]=0;ram[40][123]=0;ram[40][124]=0;ram[40][125]=0;ram[40][126]=0;ram[40][127]=0;ram[40][128]=0;ram[40][129]=0;ram[40][130]=0;ram[40][131]=0;ram[40][132]=0;ram[40][133]=0;ram[40][134]=0;ram[40][135]=0;ram[40][136]=0;ram[40][137]=0;ram[40][138]=0;ram[40][139]=0;ram[40][140]=0;
        ram[41][0]=0;ram[41][1]=0;ram[41][2]=0;ram[41][3]=0;ram[41][4]=0;ram[41][5]=0;ram[41][6]=0;ram[41][7]=0;ram[41][8]=0;ram[41][9]=0;ram[41][10]=0;ram[41][11]=0;ram[41][12]=0;ram[41][13]=0;ram[41][14]=0;ram[41][15]=0;ram[41][16]=0;ram[41][17]=0;ram[41][18]=0;ram[41][19]=0;ram[41][20]=0;ram[41][21]=0;ram[41][22]=0;ram[41][23]=0;ram[41][24]=0;ram[41][25]=0;ram[41][26]=0;ram[41][27]=0;ram[41][28]=0;ram[41][29]=1;ram[41][30]=0;ram[41][31]=0;ram[41][32]=0;ram[41][33]=0;ram[41][34]=0;ram[41][35]=1;ram[41][36]=0;ram[41][37]=1;ram[41][38]=0;ram[41][39]=1;ram[41][40]=0;ram[41][41]=1;ram[41][42]=0;ram[41][43]=0;ram[41][44]=0;ram[41][45]=1;ram[41][46]=0;ram[41][47]=1;ram[41][48]=0;ram[41][49]=1;ram[41][50]=0;ram[41][51]=0;ram[41][52]=0;ram[41][53]=1;ram[41][54]=0;ram[41][55]=0;ram[41][56]=0;ram[41][57]=1;ram[41][58]=0;ram[41][59]=1;ram[41][60]=0;ram[41][61]=1;ram[41][62]=0;ram[41][63]=1;ram[41][64]=0;ram[41][65]=1;ram[41][66]=0;ram[41][67]=0;ram[41][68]=0;ram[41][69]=1;ram[41][70]=0;ram[41][71]=1;ram[41][72]=0;ram[41][73]=1;ram[41][74]=0;ram[41][75]=1;ram[41][76]=0;ram[41][77]=1;ram[41][78]=0;ram[41][79]=1;ram[41][80]=0;ram[41][81]=1;ram[41][82]=0;ram[41][83]=1;ram[41][84]=0;ram[41][85]=0;ram[41][86]=0;ram[41][87]=1;ram[41][88]=0;ram[41][89]=0;ram[41][90]=0;ram[41][91]=1;ram[41][92]=0;ram[41][93]=1;ram[41][94]=0;ram[41][95]=0;ram[41][96]=0;ram[41][97]=1;ram[41][98]=0;ram[41][99]=1;ram[41][100]=0;ram[41][101]=0;ram[41][102]=0;ram[41][103]=1;ram[41][104]=0;ram[41][105]=1;ram[41][106]=0;ram[41][107]=1;ram[41][108]=0;ram[41][109]=1;ram[41][110]=0;ram[41][111]=1;ram[41][112]=0;ram[41][113]=0;ram[41][114]=0;ram[41][115]=0;ram[41][116]=0;ram[41][117]=0;ram[41][118]=0;ram[41][119]=0;ram[41][120]=0;ram[41][121]=0;ram[41][122]=0;ram[41][123]=0;ram[41][124]=0;ram[41][125]=0;ram[41][126]=0;ram[41][127]=0;ram[41][128]=0;ram[41][129]=0;ram[41][130]=0;ram[41][131]=0;ram[41][132]=0;ram[41][133]=0;ram[41][134]=0;ram[41][135]=0;ram[41][136]=0;ram[41][137]=0;ram[41][138]=0;ram[41][139]=0;ram[41][140]=0;
        ram[42][0]=0;ram[42][1]=0;ram[42][2]=0;ram[42][3]=0;ram[42][4]=0;ram[42][5]=0;ram[42][6]=0;ram[42][7]=0;ram[42][8]=0;ram[42][9]=0;ram[42][10]=0;ram[42][11]=0;ram[42][12]=0;ram[42][13]=0;ram[42][14]=0;ram[42][15]=0;ram[42][16]=0;ram[42][17]=0;ram[42][18]=0;ram[42][19]=0;ram[42][20]=0;ram[42][21]=0;ram[42][22]=0;ram[42][23]=0;ram[42][24]=0;ram[42][25]=0;ram[42][26]=0;ram[42][27]=0;ram[42][28]=1;ram[42][29]=0;ram[42][30]=0;ram[42][31]=0;ram[42][32]=0;ram[42][33]=0;ram[42][34]=1;ram[42][35]=0;ram[42][36]=1;ram[42][37]=0;ram[42][38]=1;ram[42][39]=0;ram[42][40]=0;ram[42][41]=0;ram[42][42]=1;ram[42][43]=0;ram[42][44]=0;ram[42][45]=0;ram[42][46]=1;ram[42][47]=0;ram[42][48]=0;ram[42][49]=0;ram[42][50]=1;ram[42][51]=0;ram[42][52]=1;ram[42][53]=0;ram[42][54]=1;ram[42][55]=0;ram[42][56]=1;ram[42][57]=0;ram[42][58]=0;ram[42][59]=0;ram[42][60]=1;ram[42][61]=0;ram[42][62]=1;ram[42][63]=0;ram[42][64]=0;ram[42][65]=0;ram[42][66]=0;ram[42][67]=0;ram[42][68]=1;ram[42][69]=0;ram[42][70]=1;ram[42][71]=0;ram[42][72]=1;ram[42][73]=0;ram[42][74]=0;ram[42][75]=0;ram[42][76]=0;ram[42][77]=0;ram[42][78]=1;ram[42][79]=0;ram[42][80]=1;ram[42][81]=0;ram[42][82]=0;ram[42][83]=0;ram[42][84]=1;ram[42][85]=0;ram[42][86]=1;ram[42][87]=0;ram[42][88]=0;ram[42][89]=0;ram[42][90]=1;ram[42][91]=0;ram[42][92]=0;ram[42][93]=0;ram[42][94]=0;ram[42][95]=0;ram[42][96]=1;ram[42][97]=0;ram[42][98]=0;ram[42][99]=0;ram[42][100]=1;ram[42][101]=0;ram[42][102]=1;ram[42][103]=0;ram[42][104]=1;ram[42][105]=0;ram[42][106]=1;ram[42][107]=0;ram[42][108]=0;ram[42][109]=0;ram[42][110]=0;ram[42][111]=0;ram[42][112]=1;ram[42][113]=0;ram[42][114]=0;ram[42][115]=0;ram[42][116]=0;ram[42][117]=0;ram[42][118]=0;ram[42][119]=0;ram[42][120]=0;ram[42][121]=0;ram[42][122]=0;ram[42][123]=0;ram[42][124]=0;ram[42][125]=0;ram[42][126]=0;ram[42][127]=0;ram[42][128]=0;ram[42][129]=0;ram[42][130]=0;ram[42][131]=0;ram[42][132]=0;ram[42][133]=0;ram[42][134]=0;ram[42][135]=0;ram[42][136]=0;ram[42][137]=0;ram[42][138]=0;ram[42][139]=0;ram[42][140]=0;
        ram[43][0]=0;ram[43][1]=0;ram[43][2]=0;ram[43][3]=0;ram[43][4]=0;ram[43][5]=0;ram[43][6]=0;ram[43][7]=0;ram[43][8]=0;ram[43][9]=0;ram[43][10]=0;ram[43][11]=0;ram[43][12]=0;ram[43][13]=0;ram[43][14]=0;ram[43][15]=0;ram[43][16]=0;ram[43][17]=0;ram[43][18]=0;ram[43][19]=0;ram[43][20]=0;ram[43][21]=0;ram[43][22]=0;ram[43][23]=0;ram[43][24]=0;ram[43][25]=0;ram[43][26]=0;ram[43][27]=1;ram[43][28]=0;ram[43][29]=1;ram[43][30]=0;ram[43][31]=0;ram[43][32]=0;ram[43][33]=1;ram[43][34]=0;ram[43][35]=0;ram[43][36]=0;ram[43][37]=1;ram[43][38]=0;ram[43][39]=1;ram[43][40]=0;ram[43][41]=1;ram[43][42]=0;ram[43][43]=1;ram[43][44]=0;ram[43][45]=0;ram[43][46]=0;ram[43][47]=1;ram[43][48]=0;ram[43][49]=0;ram[43][50]=0;ram[43][51]=1;ram[43][52]=0;ram[43][53]=1;ram[43][54]=0;ram[43][55]=0;ram[43][56]=0;ram[43][57]=1;ram[43][58]=0;ram[43][59]=1;ram[43][60]=0;ram[43][61]=1;ram[43][62]=0;ram[43][63]=0;ram[43][64]=0;ram[43][65]=1;ram[43][66]=0;ram[43][67]=1;ram[43][68]=0;ram[43][69]=1;ram[43][70]=0;ram[43][71]=0;ram[43][72]=0;ram[43][73]=1;ram[43][74]=0;ram[43][75]=1;ram[43][76]=0;ram[43][77]=1;ram[43][78]=0;ram[43][79]=0;ram[43][80]=0;ram[43][81]=0;ram[43][82]=0;ram[43][83]=1;ram[43][84]=0;ram[43][85]=1;ram[43][86]=0;ram[43][87]=1;ram[43][88]=0;ram[43][89]=1;ram[43][90]=0;ram[43][91]=1;ram[43][92]=0;ram[43][93]=1;ram[43][94]=0;ram[43][95]=0;ram[43][96]=0;ram[43][97]=1;ram[43][98]=0;ram[43][99]=1;ram[43][100]=0;ram[43][101]=0;ram[43][102]=0;ram[43][103]=0;ram[43][104]=0;ram[43][105]=1;ram[43][106]=0;ram[43][107]=1;ram[43][108]=0;ram[43][109]=1;ram[43][110]=0;ram[43][111]=0;ram[43][112]=0;ram[43][113]=1;ram[43][114]=0;ram[43][115]=0;ram[43][116]=0;ram[43][117]=0;ram[43][118]=0;ram[43][119]=0;ram[43][120]=0;ram[43][121]=0;ram[43][122]=0;ram[43][123]=0;ram[43][124]=0;ram[43][125]=0;ram[43][126]=0;ram[43][127]=0;ram[43][128]=0;ram[43][129]=0;ram[43][130]=0;ram[43][131]=0;ram[43][132]=0;ram[43][133]=0;ram[43][134]=0;ram[43][135]=0;ram[43][136]=0;ram[43][137]=0;ram[43][138]=0;ram[43][139]=0;ram[43][140]=0;
        ram[44][0]=0;ram[44][1]=0;ram[44][2]=0;ram[44][3]=0;ram[44][4]=0;ram[44][5]=0;ram[44][6]=0;ram[44][7]=0;ram[44][8]=0;ram[44][9]=0;ram[44][10]=0;ram[44][11]=0;ram[44][12]=0;ram[44][13]=0;ram[44][14]=0;ram[44][15]=0;ram[44][16]=0;ram[44][17]=0;ram[44][18]=0;ram[44][19]=0;ram[44][20]=0;ram[44][21]=0;ram[44][22]=0;ram[44][23]=0;ram[44][24]=0;ram[44][25]=0;ram[44][26]=1;ram[44][27]=0;ram[44][28]=0;ram[44][29]=0;ram[44][30]=1;ram[44][31]=0;ram[44][32]=0;ram[44][33]=0;ram[44][34]=0;ram[44][35]=0;ram[44][36]=1;ram[44][37]=0;ram[44][38]=0;ram[44][39]=0;ram[44][40]=1;ram[44][41]=0;ram[44][42]=1;ram[44][43]=0;ram[44][44]=1;ram[44][45]=0;ram[44][46]=0;ram[44][47]=0;ram[44][48]=1;ram[44][49]=0;ram[44][50]=0;ram[44][51]=0;ram[44][52]=1;ram[44][53]=0;ram[44][54]=1;ram[44][55]=0;ram[44][56]=1;ram[44][57]=0;ram[44][58]=1;ram[44][59]=0;ram[44][60]=1;ram[44][61]=0;ram[44][62]=1;ram[44][63]=0;ram[44][64]=0;ram[44][65]=0;ram[44][66]=1;ram[44][67]=0;ram[44][68]=1;ram[44][69]=0;ram[44][70]=1;ram[44][71]=0;ram[44][72]=0;ram[44][73]=0;ram[44][74]=1;ram[44][75]=0;ram[44][76]=1;ram[44][77]=0;ram[44][78]=0;ram[44][79]=0;ram[44][80]=1;ram[44][81]=0;ram[44][82]=0;ram[44][83]=0;ram[44][84]=0;ram[44][85]=0;ram[44][86]=1;ram[44][87]=0;ram[44][88]=0;ram[44][89]=0;ram[44][90]=1;ram[44][91]=0;ram[44][92]=1;ram[44][93]=0;ram[44][94]=1;ram[44][95]=0;ram[44][96]=1;ram[44][97]=0;ram[44][98]=1;ram[44][99]=0;ram[44][100]=1;ram[44][101]=0;ram[44][102]=1;ram[44][103]=0;ram[44][104]=1;ram[44][105]=0;ram[44][106]=1;ram[44][107]=0;ram[44][108]=1;ram[44][109]=0;ram[44][110]=1;ram[44][111]=0;ram[44][112]=1;ram[44][113]=0;ram[44][114]=1;ram[44][115]=0;ram[44][116]=0;ram[44][117]=0;ram[44][118]=0;ram[44][119]=0;ram[44][120]=0;ram[44][121]=0;ram[44][122]=0;ram[44][123]=0;ram[44][124]=0;ram[44][125]=0;ram[44][126]=0;ram[44][127]=0;ram[44][128]=0;ram[44][129]=0;ram[44][130]=0;ram[44][131]=0;ram[44][132]=0;ram[44][133]=0;ram[44][134]=0;ram[44][135]=0;ram[44][136]=0;ram[44][137]=0;ram[44][138]=0;ram[44][139]=0;ram[44][140]=0;
        ram[45][0]=0;ram[45][1]=0;ram[45][2]=0;ram[45][3]=0;ram[45][4]=0;ram[45][5]=0;ram[45][6]=0;ram[45][7]=0;ram[45][8]=0;ram[45][9]=0;ram[45][10]=0;ram[45][11]=0;ram[45][12]=0;ram[45][13]=0;ram[45][14]=0;ram[45][15]=0;ram[45][16]=0;ram[45][17]=0;ram[45][18]=0;ram[45][19]=0;ram[45][20]=0;ram[45][21]=0;ram[45][22]=0;ram[45][23]=0;ram[45][24]=0;ram[45][25]=1;ram[45][26]=0;ram[45][27]=1;ram[45][28]=0;ram[45][29]=0;ram[45][30]=0;ram[45][31]=0;ram[45][32]=0;ram[45][33]=1;ram[45][34]=0;ram[45][35]=1;ram[45][36]=0;ram[45][37]=1;ram[45][38]=0;ram[45][39]=0;ram[45][40]=0;ram[45][41]=0;ram[45][42]=0;ram[45][43]=1;ram[45][44]=0;ram[45][45]=1;ram[45][46]=0;ram[45][47]=1;ram[45][48]=0;ram[45][49]=1;ram[45][50]=0;ram[45][51]=1;ram[45][52]=0;ram[45][53]=1;ram[45][54]=0;ram[45][55]=1;ram[45][56]=0;ram[45][57]=1;ram[45][58]=0;ram[45][59]=0;ram[45][60]=0;ram[45][61]=1;ram[45][62]=0;ram[45][63]=0;ram[45][64]=0;ram[45][65]=1;ram[45][66]=0;ram[45][67]=1;ram[45][68]=0;ram[45][69]=0;ram[45][70]=0;ram[45][71]=0;ram[45][72]=0;ram[45][73]=1;ram[45][74]=0;ram[45][75]=0;ram[45][76]=0;ram[45][77]=1;ram[45][78]=0;ram[45][79]=1;ram[45][80]=0;ram[45][81]=1;ram[45][82]=0;ram[45][83]=0;ram[45][84]=0;ram[45][85]=0;ram[45][86]=0;ram[45][87]=1;ram[45][88]=0;ram[45][89]=1;ram[45][90]=0;ram[45][91]=1;ram[45][92]=0;ram[45][93]=0;ram[45][94]=0;ram[45][95]=1;ram[45][96]=0;ram[45][97]=1;ram[45][98]=0;ram[45][99]=1;ram[45][100]=0;ram[45][101]=0;ram[45][102]=0;ram[45][103]=1;ram[45][104]=0;ram[45][105]=1;ram[45][106]=0;ram[45][107]=0;ram[45][108]=0;ram[45][109]=1;ram[45][110]=0;ram[45][111]=1;ram[45][112]=0;ram[45][113]=0;ram[45][114]=0;ram[45][115]=1;ram[45][116]=0;ram[45][117]=0;ram[45][118]=0;ram[45][119]=0;ram[45][120]=0;ram[45][121]=0;ram[45][122]=0;ram[45][123]=0;ram[45][124]=0;ram[45][125]=0;ram[45][126]=0;ram[45][127]=0;ram[45][128]=0;ram[45][129]=0;ram[45][130]=0;ram[45][131]=0;ram[45][132]=0;ram[45][133]=0;ram[45][134]=0;ram[45][135]=0;ram[45][136]=0;ram[45][137]=0;ram[45][138]=0;ram[45][139]=0;ram[45][140]=0;
        ram[46][0]=0;ram[46][1]=0;ram[46][2]=0;ram[46][3]=0;ram[46][4]=0;ram[46][5]=0;ram[46][6]=0;ram[46][7]=0;ram[46][8]=0;ram[46][9]=0;ram[46][10]=0;ram[46][11]=0;ram[46][12]=0;ram[46][13]=0;ram[46][14]=0;ram[46][15]=0;ram[46][16]=0;ram[46][17]=0;ram[46][18]=0;ram[46][19]=0;ram[46][20]=0;ram[46][21]=0;ram[46][22]=0;ram[46][23]=0;ram[46][24]=1;ram[46][25]=0;ram[46][26]=1;ram[46][27]=0;ram[46][28]=1;ram[46][29]=0;ram[46][30]=0;ram[46][31]=0;ram[46][32]=1;ram[46][33]=0;ram[46][34]=1;ram[46][35]=0;ram[46][36]=1;ram[46][37]=0;ram[46][38]=1;ram[46][39]=0;ram[46][40]=1;ram[46][41]=0;ram[46][42]=1;ram[46][43]=0;ram[46][44]=1;ram[46][45]=0;ram[46][46]=1;ram[46][47]=0;ram[46][48]=1;ram[46][49]=0;ram[46][50]=0;ram[46][51]=0;ram[46][52]=1;ram[46][53]=0;ram[46][54]=0;ram[46][55]=0;ram[46][56]=1;ram[46][57]=0;ram[46][58]=1;ram[46][59]=0;ram[46][60]=1;ram[46][61]=0;ram[46][62]=1;ram[46][63]=0;ram[46][64]=1;ram[46][65]=0;ram[46][66]=1;ram[46][67]=0;ram[46][68]=0;ram[46][69]=0;ram[46][70]=1;ram[46][71]=0;ram[46][72]=1;ram[46][73]=0;ram[46][74]=0;ram[46][75]=0;ram[46][76]=1;ram[46][77]=0;ram[46][78]=1;ram[46][79]=0;ram[46][80]=1;ram[46][81]=0;ram[46][82]=1;ram[46][83]=0;ram[46][84]=0;ram[46][85]=0;ram[46][86]=0;ram[46][87]=0;ram[46][88]=1;ram[46][89]=0;ram[46][90]=1;ram[46][91]=0;ram[46][92]=1;ram[46][93]=0;ram[46][94]=1;ram[46][95]=0;ram[46][96]=1;ram[46][97]=0;ram[46][98]=0;ram[46][99]=0;ram[46][100]=1;ram[46][101]=0;ram[46][102]=0;ram[46][103]=0;ram[46][104]=1;ram[46][105]=0;ram[46][106]=0;ram[46][107]=0;ram[46][108]=1;ram[46][109]=0;ram[46][110]=1;ram[46][111]=0;ram[46][112]=0;ram[46][113]=0;ram[46][114]=0;ram[46][115]=0;ram[46][116]=1;ram[46][117]=0;ram[46][118]=0;ram[46][119]=0;ram[46][120]=0;ram[46][121]=0;ram[46][122]=0;ram[46][123]=0;ram[46][124]=0;ram[46][125]=0;ram[46][126]=0;ram[46][127]=0;ram[46][128]=0;ram[46][129]=0;ram[46][130]=0;ram[46][131]=0;ram[46][132]=0;ram[46][133]=0;ram[46][134]=0;ram[46][135]=0;ram[46][136]=0;ram[46][137]=0;ram[46][138]=0;ram[46][139]=0;ram[46][140]=0;
        ram[47][0]=0;ram[47][1]=0;ram[47][2]=0;ram[47][3]=0;ram[47][4]=0;ram[47][5]=0;ram[47][6]=0;ram[47][7]=0;ram[47][8]=0;ram[47][9]=0;ram[47][10]=0;ram[47][11]=0;ram[47][12]=0;ram[47][13]=0;ram[47][14]=0;ram[47][15]=0;ram[47][16]=0;ram[47][17]=0;ram[47][18]=0;ram[47][19]=0;ram[47][20]=0;ram[47][21]=0;ram[47][22]=0;ram[47][23]=1;ram[47][24]=0;ram[47][25]=1;ram[47][26]=0;ram[47][27]=0;ram[47][28]=0;ram[47][29]=1;ram[47][30]=0;ram[47][31]=1;ram[47][32]=0;ram[47][33]=1;ram[47][34]=0;ram[47][35]=0;ram[47][36]=0;ram[47][37]=1;ram[47][38]=0;ram[47][39]=0;ram[47][40]=0;ram[47][41]=1;ram[47][42]=0;ram[47][43]=0;ram[47][44]=0;ram[47][45]=1;ram[47][46]=0;ram[47][47]=1;ram[47][48]=0;ram[47][49]=1;ram[47][50]=0;ram[47][51]=1;ram[47][52]=0;ram[47][53]=0;ram[47][54]=0;ram[47][55]=0;ram[47][56]=0;ram[47][57]=1;ram[47][58]=0;ram[47][59]=1;ram[47][60]=0;ram[47][61]=1;ram[47][62]=0;ram[47][63]=0;ram[47][64]=0;ram[47][65]=1;ram[47][66]=0;ram[47][67]=0;ram[47][68]=0;ram[47][69]=0;ram[47][70]=0;ram[47][71]=1;ram[47][72]=0;ram[47][73]=0;ram[47][74]=0;ram[47][75]=1;ram[47][76]=0;ram[47][77]=1;ram[47][78]=0;ram[47][79]=1;ram[47][80]=0;ram[47][81]=1;ram[47][82]=0;ram[47][83]=0;ram[47][84]=0;ram[47][85]=1;ram[47][86]=0;ram[47][87]=0;ram[47][88]=0;ram[47][89]=1;ram[47][90]=0;ram[47][91]=1;ram[47][92]=0;ram[47][93]=0;ram[47][94]=0;ram[47][95]=0;ram[47][96]=0;ram[47][97]=1;ram[47][98]=0;ram[47][99]=1;ram[47][100]=0;ram[47][101]=1;ram[47][102]=0;ram[47][103]=1;ram[47][104]=0;ram[47][105]=1;ram[47][106]=0;ram[47][107]=1;ram[47][108]=0;ram[47][109]=1;ram[47][110]=0;ram[47][111]=1;ram[47][112]=0;ram[47][113]=0;ram[47][114]=0;ram[47][115]=1;ram[47][116]=0;ram[47][117]=1;ram[47][118]=0;ram[47][119]=0;ram[47][120]=0;ram[47][121]=0;ram[47][122]=0;ram[47][123]=0;ram[47][124]=0;ram[47][125]=0;ram[47][126]=0;ram[47][127]=0;ram[47][128]=0;ram[47][129]=0;ram[47][130]=0;ram[47][131]=0;ram[47][132]=0;ram[47][133]=0;ram[47][134]=0;ram[47][135]=0;ram[47][136]=0;ram[47][137]=0;ram[47][138]=0;ram[47][139]=0;ram[47][140]=0;
        ram[48][0]=0;ram[48][1]=0;ram[48][2]=0;ram[48][3]=0;ram[48][4]=0;ram[48][5]=0;ram[48][6]=0;ram[48][7]=0;ram[48][8]=0;ram[48][9]=0;ram[48][10]=0;ram[48][11]=0;ram[48][12]=0;ram[48][13]=0;ram[48][14]=0;ram[48][15]=0;ram[48][16]=0;ram[48][17]=0;ram[48][18]=0;ram[48][19]=0;ram[48][20]=0;ram[48][21]=0;ram[48][22]=1;ram[48][23]=0;ram[48][24]=1;ram[48][25]=0;ram[48][26]=1;ram[48][27]=0;ram[48][28]=1;ram[48][29]=0;ram[48][30]=1;ram[48][31]=0;ram[48][32]=0;ram[48][33]=0;ram[48][34]=1;ram[48][35]=0;ram[48][36]=0;ram[48][37]=0;ram[48][38]=1;ram[48][39]=0;ram[48][40]=1;ram[48][41]=0;ram[48][42]=1;ram[48][43]=0;ram[48][44]=0;ram[48][45]=0;ram[48][46]=1;ram[48][47]=0;ram[48][48]=1;ram[48][49]=0;ram[48][50]=1;ram[48][51]=0;ram[48][52]=0;ram[48][53]=0;ram[48][54]=1;ram[48][55]=0;ram[48][56]=0;ram[48][57]=0;ram[48][58]=1;ram[48][59]=0;ram[48][60]=1;ram[48][61]=0;ram[48][62]=0;ram[48][63]=0;ram[48][64]=0;ram[48][65]=0;ram[48][66]=1;ram[48][67]=0;ram[48][68]=1;ram[48][69]=0;ram[48][70]=0;ram[48][71]=0;ram[48][72]=0;ram[48][73]=0;ram[48][74]=1;ram[48][75]=0;ram[48][76]=1;ram[48][77]=0;ram[48][78]=1;ram[48][79]=0;ram[48][80]=1;ram[48][81]=0;ram[48][82]=0;ram[48][83]=0;ram[48][84]=1;ram[48][85]=0;ram[48][86]=1;ram[48][87]=0;ram[48][88]=1;ram[48][89]=0;ram[48][90]=1;ram[48][91]=0;ram[48][92]=1;ram[48][93]=0;ram[48][94]=1;ram[48][95]=0;ram[48][96]=0;ram[48][97]=0;ram[48][98]=1;ram[48][99]=0;ram[48][100]=1;ram[48][101]=0;ram[48][102]=0;ram[48][103]=0;ram[48][104]=1;ram[48][105]=0;ram[48][106]=0;ram[48][107]=0;ram[48][108]=1;ram[48][109]=0;ram[48][110]=1;ram[48][111]=0;ram[48][112]=0;ram[48][113]=0;ram[48][114]=0;ram[48][115]=0;ram[48][116]=1;ram[48][117]=0;ram[48][118]=1;ram[48][119]=0;ram[48][120]=0;ram[48][121]=0;ram[48][122]=0;ram[48][123]=0;ram[48][124]=0;ram[48][125]=0;ram[48][126]=0;ram[48][127]=0;ram[48][128]=0;ram[48][129]=0;ram[48][130]=0;ram[48][131]=0;ram[48][132]=0;ram[48][133]=0;ram[48][134]=0;ram[48][135]=0;ram[48][136]=0;ram[48][137]=0;ram[48][138]=0;ram[48][139]=0;ram[48][140]=0;
        ram[49][0]=0;ram[49][1]=0;ram[49][2]=0;ram[49][3]=0;ram[49][4]=0;ram[49][5]=0;ram[49][6]=0;ram[49][7]=0;ram[49][8]=0;ram[49][9]=0;ram[49][10]=0;ram[49][11]=0;ram[49][12]=0;ram[49][13]=0;ram[49][14]=0;ram[49][15]=0;ram[49][16]=0;ram[49][17]=0;ram[49][18]=0;ram[49][19]=0;ram[49][20]=0;ram[49][21]=1;ram[49][22]=0;ram[49][23]=0;ram[49][24]=0;ram[49][25]=1;ram[49][26]=0;ram[49][27]=0;ram[49][28]=0;ram[49][29]=0;ram[49][30]=0;ram[49][31]=1;ram[49][32]=0;ram[49][33]=0;ram[49][34]=0;ram[49][35]=1;ram[49][36]=0;ram[49][37]=0;ram[49][38]=0;ram[49][39]=1;ram[49][40]=0;ram[49][41]=1;ram[49][42]=0;ram[49][43]=0;ram[49][44]=0;ram[49][45]=1;ram[49][46]=0;ram[49][47]=1;ram[49][48]=0;ram[49][49]=1;ram[49][50]=0;ram[49][51]=1;ram[49][52]=0;ram[49][53]=1;ram[49][54]=0;ram[49][55]=0;ram[49][56]=0;ram[49][57]=0;ram[49][58]=0;ram[49][59]=1;ram[49][60]=0;ram[49][61]=1;ram[49][62]=0;ram[49][63]=1;ram[49][64]=0;ram[49][65]=1;ram[49][66]=0;ram[49][67]=1;ram[49][68]=0;ram[49][69]=1;ram[49][70]=0;ram[49][71]=1;ram[49][72]=0;ram[49][73]=1;ram[49][74]=0;ram[49][75]=1;ram[49][76]=0;ram[49][77]=1;ram[49][78]=0;ram[49][79]=1;ram[49][80]=0;ram[49][81]=1;ram[49][82]=0;ram[49][83]=1;ram[49][84]=0;ram[49][85]=1;ram[49][86]=0;ram[49][87]=0;ram[49][88]=0;ram[49][89]=0;ram[49][90]=0;ram[49][91]=1;ram[49][92]=0;ram[49][93]=1;ram[49][94]=0;ram[49][95]=1;ram[49][96]=0;ram[49][97]=1;ram[49][98]=0;ram[49][99]=1;ram[49][100]=0;ram[49][101]=1;ram[49][102]=0;ram[49][103]=1;ram[49][104]=0;ram[49][105]=1;ram[49][106]=0;ram[49][107]=1;ram[49][108]=0;ram[49][109]=0;ram[49][110]=0;ram[49][111]=0;ram[49][112]=0;ram[49][113]=0;ram[49][114]=0;ram[49][115]=1;ram[49][116]=0;ram[49][117]=0;ram[49][118]=0;ram[49][119]=1;ram[49][120]=0;ram[49][121]=0;ram[49][122]=0;ram[49][123]=0;ram[49][124]=0;ram[49][125]=0;ram[49][126]=0;ram[49][127]=0;ram[49][128]=0;ram[49][129]=0;ram[49][130]=0;ram[49][131]=0;ram[49][132]=0;ram[49][133]=0;ram[49][134]=0;ram[49][135]=0;ram[49][136]=0;ram[49][137]=0;ram[49][138]=0;ram[49][139]=0;ram[49][140]=0;
        ram[50][0]=0;ram[50][1]=0;ram[50][2]=0;ram[50][3]=0;ram[50][4]=0;ram[50][5]=0;ram[50][6]=0;ram[50][7]=0;ram[50][8]=0;ram[50][9]=0;ram[50][10]=0;ram[50][11]=0;ram[50][12]=0;ram[50][13]=0;ram[50][14]=0;ram[50][15]=0;ram[50][16]=0;ram[50][17]=0;ram[50][18]=0;ram[50][19]=0;ram[50][20]=1;ram[50][21]=0;ram[50][22]=1;ram[50][23]=0;ram[50][24]=1;ram[50][25]=0;ram[50][26]=0;ram[50][27]=0;ram[50][28]=0;ram[50][29]=0;ram[50][30]=1;ram[50][31]=0;ram[50][32]=1;ram[50][33]=0;ram[50][34]=1;ram[50][35]=0;ram[50][36]=0;ram[50][37]=0;ram[50][38]=1;ram[50][39]=0;ram[50][40]=1;ram[50][41]=0;ram[50][42]=0;ram[50][43]=0;ram[50][44]=1;ram[50][45]=0;ram[50][46]=1;ram[50][47]=0;ram[50][48]=1;ram[50][49]=0;ram[50][50]=1;ram[50][51]=0;ram[50][52]=1;ram[50][53]=0;ram[50][54]=0;ram[50][55]=0;ram[50][56]=0;ram[50][57]=0;ram[50][58]=1;ram[50][59]=0;ram[50][60]=0;ram[50][61]=0;ram[50][62]=1;ram[50][63]=0;ram[50][64]=0;ram[50][65]=0;ram[50][66]=1;ram[50][67]=0;ram[50][68]=1;ram[50][69]=0;ram[50][70]=0;ram[50][71]=0;ram[50][72]=0;ram[50][73]=0;ram[50][74]=1;ram[50][75]=0;ram[50][76]=1;ram[50][77]=0;ram[50][78]=1;ram[50][79]=0;ram[50][80]=1;ram[50][81]=0;ram[50][82]=0;ram[50][83]=0;ram[50][84]=1;ram[50][85]=0;ram[50][86]=1;ram[50][87]=0;ram[50][88]=0;ram[50][89]=0;ram[50][90]=1;ram[50][91]=0;ram[50][92]=0;ram[50][93]=0;ram[50][94]=1;ram[50][95]=0;ram[50][96]=0;ram[50][97]=0;ram[50][98]=1;ram[50][99]=0;ram[50][100]=1;ram[50][101]=0;ram[50][102]=1;ram[50][103]=0;ram[50][104]=1;ram[50][105]=0;ram[50][106]=1;ram[50][107]=0;ram[50][108]=0;ram[50][109]=0;ram[50][110]=1;ram[50][111]=0;ram[50][112]=0;ram[50][113]=0;ram[50][114]=0;ram[50][115]=0;ram[50][116]=0;ram[50][117]=0;ram[50][118]=1;ram[50][119]=0;ram[50][120]=1;ram[50][121]=0;ram[50][122]=0;ram[50][123]=0;ram[50][124]=0;ram[50][125]=0;ram[50][126]=0;ram[50][127]=0;ram[50][128]=0;ram[50][129]=0;ram[50][130]=0;ram[50][131]=0;ram[50][132]=0;ram[50][133]=0;ram[50][134]=0;ram[50][135]=0;ram[50][136]=0;ram[50][137]=0;ram[50][138]=0;ram[50][139]=0;ram[50][140]=0;
        ram[51][0]=0;ram[51][1]=0;ram[51][2]=0;ram[51][3]=0;ram[51][4]=0;ram[51][5]=0;ram[51][6]=0;ram[51][7]=0;ram[51][8]=0;ram[51][9]=0;ram[51][10]=0;ram[51][11]=0;ram[51][12]=0;ram[51][13]=0;ram[51][14]=0;ram[51][15]=0;ram[51][16]=0;ram[51][17]=0;ram[51][18]=0;ram[51][19]=1;ram[51][20]=0;ram[51][21]=0;ram[51][22]=0;ram[51][23]=1;ram[51][24]=0;ram[51][25]=1;ram[51][26]=0;ram[51][27]=1;ram[51][28]=0;ram[51][29]=1;ram[51][30]=0;ram[51][31]=1;ram[51][32]=0;ram[51][33]=1;ram[51][34]=0;ram[51][35]=0;ram[51][36]=0;ram[51][37]=1;ram[51][38]=0;ram[51][39]=1;ram[51][40]=0;ram[51][41]=1;ram[51][42]=0;ram[51][43]=0;ram[51][44]=0;ram[51][45]=1;ram[51][46]=0;ram[51][47]=0;ram[51][48]=0;ram[51][49]=1;ram[51][50]=0;ram[51][51]=1;ram[51][52]=0;ram[51][53]=1;ram[51][54]=0;ram[51][55]=1;ram[51][56]=0;ram[51][57]=1;ram[51][58]=0;ram[51][59]=1;ram[51][60]=0;ram[51][61]=0;ram[51][62]=0;ram[51][63]=0;ram[51][64]=0;ram[51][65]=1;ram[51][66]=0;ram[51][67]=1;ram[51][68]=0;ram[51][69]=0;ram[51][70]=0;ram[51][71]=0;ram[51][72]=0;ram[51][73]=0;ram[51][74]=0;ram[51][75]=1;ram[51][76]=0;ram[51][77]=0;ram[51][78]=0;ram[51][79]=0;ram[51][80]=0;ram[51][81]=1;ram[51][82]=0;ram[51][83]=0;ram[51][84]=0;ram[51][85]=1;ram[51][86]=0;ram[51][87]=1;ram[51][88]=0;ram[51][89]=0;ram[51][90]=0;ram[51][91]=1;ram[51][92]=0;ram[51][93]=1;ram[51][94]=0;ram[51][95]=0;ram[51][96]=0;ram[51][97]=1;ram[51][98]=0;ram[51][99]=0;ram[51][100]=0;ram[51][101]=1;ram[51][102]=0;ram[51][103]=1;ram[51][104]=0;ram[51][105]=1;ram[51][106]=0;ram[51][107]=1;ram[51][108]=0;ram[51][109]=1;ram[51][110]=0;ram[51][111]=0;ram[51][112]=0;ram[51][113]=1;ram[51][114]=0;ram[51][115]=1;ram[51][116]=0;ram[51][117]=0;ram[51][118]=0;ram[51][119]=1;ram[51][120]=0;ram[51][121]=1;ram[51][122]=0;ram[51][123]=0;ram[51][124]=0;ram[51][125]=0;ram[51][126]=0;ram[51][127]=0;ram[51][128]=0;ram[51][129]=0;ram[51][130]=0;ram[51][131]=0;ram[51][132]=0;ram[51][133]=0;ram[51][134]=0;ram[51][135]=0;ram[51][136]=0;ram[51][137]=0;ram[51][138]=0;ram[51][139]=0;ram[51][140]=0;
        ram[52][0]=0;ram[52][1]=0;ram[52][2]=0;ram[52][3]=0;ram[52][4]=0;ram[52][5]=0;ram[52][6]=0;ram[52][7]=0;ram[52][8]=0;ram[52][9]=0;ram[52][10]=0;ram[52][11]=0;ram[52][12]=0;ram[52][13]=0;ram[52][14]=0;ram[52][15]=0;ram[52][16]=0;ram[52][17]=0;ram[52][18]=1;ram[52][19]=0;ram[52][20]=1;ram[52][21]=0;ram[52][22]=1;ram[52][23]=0;ram[52][24]=1;ram[52][25]=0;ram[52][26]=1;ram[52][27]=0;ram[52][28]=1;ram[52][29]=0;ram[52][30]=1;ram[52][31]=0;ram[52][32]=1;ram[52][33]=0;ram[52][34]=1;ram[52][35]=0;ram[52][36]=0;ram[52][37]=0;ram[52][38]=0;ram[52][39]=0;ram[52][40]=1;ram[52][41]=0;ram[52][42]=0;ram[52][43]=0;ram[52][44]=0;ram[52][45]=0;ram[52][46]=0;ram[52][47]=0;ram[52][48]=0;ram[52][49]=0;ram[52][50]=1;ram[52][51]=0;ram[52][52]=1;ram[52][53]=0;ram[52][54]=0;ram[52][55]=0;ram[52][56]=0;ram[52][57]=0;ram[52][58]=1;ram[52][59]=0;ram[52][60]=1;ram[52][61]=0;ram[52][62]=1;ram[52][63]=0;ram[52][64]=1;ram[52][65]=0;ram[52][66]=1;ram[52][67]=0;ram[52][68]=1;ram[52][69]=0;ram[52][70]=1;ram[52][71]=0;ram[52][72]=1;ram[52][73]=0;ram[52][74]=0;ram[52][75]=0;ram[52][76]=1;ram[52][77]=0;ram[52][78]=0;ram[52][79]=0;ram[52][80]=1;ram[52][81]=0;ram[52][82]=1;ram[52][83]=0;ram[52][84]=0;ram[52][85]=0;ram[52][86]=1;ram[52][87]=0;ram[52][88]=0;ram[52][89]=0;ram[52][90]=1;ram[52][91]=0;ram[52][92]=0;ram[52][93]=0;ram[52][94]=1;ram[52][95]=0;ram[52][96]=0;ram[52][97]=0;ram[52][98]=1;ram[52][99]=0;ram[52][100]=0;ram[52][101]=0;ram[52][102]=0;ram[52][103]=0;ram[52][104]=0;ram[52][105]=0;ram[52][106]=1;ram[52][107]=0;ram[52][108]=0;ram[52][109]=0;ram[52][110]=1;ram[52][111]=0;ram[52][112]=1;ram[52][113]=0;ram[52][114]=1;ram[52][115]=0;ram[52][116]=0;ram[52][117]=0;ram[52][118]=1;ram[52][119]=0;ram[52][120]=0;ram[52][121]=0;ram[52][122]=1;ram[52][123]=0;ram[52][124]=0;ram[52][125]=0;ram[52][126]=0;ram[52][127]=0;ram[52][128]=0;ram[52][129]=0;ram[52][130]=0;ram[52][131]=0;ram[52][132]=0;ram[52][133]=0;ram[52][134]=0;ram[52][135]=0;ram[52][136]=0;ram[52][137]=0;ram[52][138]=0;ram[52][139]=0;ram[52][140]=0;
        ram[53][0]=0;ram[53][1]=0;ram[53][2]=0;ram[53][3]=0;ram[53][4]=0;ram[53][5]=0;ram[53][6]=0;ram[53][7]=0;ram[53][8]=0;ram[53][9]=0;ram[53][10]=0;ram[53][11]=0;ram[53][12]=0;ram[53][13]=0;ram[53][14]=0;ram[53][15]=0;ram[53][16]=0;ram[53][17]=1;ram[53][18]=0;ram[53][19]=1;ram[53][20]=0;ram[53][21]=1;ram[53][22]=0;ram[53][23]=1;ram[53][24]=0;ram[53][25]=0;ram[53][26]=0;ram[53][27]=1;ram[53][28]=0;ram[53][29]=1;ram[53][30]=0;ram[53][31]=1;ram[53][32]=0;ram[53][33]=1;ram[53][34]=0;ram[53][35]=0;ram[53][36]=0;ram[53][37]=0;ram[53][38]=0;ram[53][39]=0;ram[53][40]=0;ram[53][41]=1;ram[53][42]=0;ram[53][43]=1;ram[53][44]=0;ram[53][45]=0;ram[53][46]=0;ram[53][47]=1;ram[53][48]=0;ram[53][49]=1;ram[53][50]=0;ram[53][51]=1;ram[53][52]=0;ram[53][53]=1;ram[53][54]=0;ram[53][55]=1;ram[53][56]=0;ram[53][57]=0;ram[53][58]=0;ram[53][59]=1;ram[53][60]=0;ram[53][61]=0;ram[53][62]=0;ram[53][63]=1;ram[53][64]=0;ram[53][65]=1;ram[53][66]=0;ram[53][67]=0;ram[53][68]=0;ram[53][69]=1;ram[53][70]=0;ram[53][71]=0;ram[53][72]=0;ram[53][73]=0;ram[53][74]=0;ram[53][75]=1;ram[53][76]=0;ram[53][77]=1;ram[53][78]=0;ram[53][79]=0;ram[53][80]=0;ram[53][81]=1;ram[53][82]=0;ram[53][83]=1;ram[53][84]=0;ram[53][85]=1;ram[53][86]=0;ram[53][87]=1;ram[53][88]=0;ram[53][89]=0;ram[53][90]=0;ram[53][91]=0;ram[53][92]=0;ram[53][93]=1;ram[53][94]=0;ram[53][95]=1;ram[53][96]=0;ram[53][97]=1;ram[53][98]=0;ram[53][99]=0;ram[53][100]=0;ram[53][101]=0;ram[53][102]=0;ram[53][103]=1;ram[53][104]=0;ram[53][105]=1;ram[53][106]=0;ram[53][107]=0;ram[53][108]=0;ram[53][109]=0;ram[53][110]=0;ram[53][111]=0;ram[53][112]=0;ram[53][113]=1;ram[53][114]=0;ram[53][115]=1;ram[53][116]=0;ram[53][117]=1;ram[53][118]=0;ram[53][119]=1;ram[53][120]=0;ram[53][121]=1;ram[53][122]=0;ram[53][123]=1;ram[53][124]=0;ram[53][125]=0;ram[53][126]=0;ram[53][127]=0;ram[53][128]=0;ram[53][129]=0;ram[53][130]=0;ram[53][131]=0;ram[53][132]=0;ram[53][133]=0;ram[53][134]=0;ram[53][135]=0;ram[53][136]=0;ram[53][137]=0;ram[53][138]=0;ram[53][139]=0;ram[53][140]=0;
        ram[54][0]=0;ram[54][1]=0;ram[54][2]=0;ram[54][3]=0;ram[54][4]=0;ram[54][5]=0;ram[54][6]=0;ram[54][7]=0;ram[54][8]=0;ram[54][9]=0;ram[54][10]=0;ram[54][11]=0;ram[54][12]=0;ram[54][13]=0;ram[54][14]=0;ram[54][15]=0;ram[54][16]=1;ram[54][17]=0;ram[54][18]=1;ram[54][19]=0;ram[54][20]=1;ram[54][21]=0;ram[54][22]=0;ram[54][23]=0;ram[54][24]=0;ram[54][25]=0;ram[54][26]=0;ram[54][27]=0;ram[54][28]=0;ram[54][29]=0;ram[54][30]=0;ram[54][31]=0;ram[54][32]=1;ram[54][33]=0;ram[54][34]=0;ram[54][35]=0;ram[54][36]=0;ram[54][37]=0;ram[54][38]=0;ram[54][39]=0;ram[54][40]=1;ram[54][41]=0;ram[54][42]=1;ram[54][43]=0;ram[54][44]=1;ram[54][45]=0;ram[54][46]=1;ram[54][47]=0;ram[54][48]=0;ram[54][49]=0;ram[54][50]=1;ram[54][51]=0;ram[54][52]=1;ram[54][53]=0;ram[54][54]=1;ram[54][55]=0;ram[54][56]=0;ram[54][57]=0;ram[54][58]=1;ram[54][59]=0;ram[54][60]=0;ram[54][61]=0;ram[54][62]=0;ram[54][63]=0;ram[54][64]=0;ram[54][65]=0;ram[54][66]=1;ram[54][67]=0;ram[54][68]=1;ram[54][69]=0;ram[54][70]=0;ram[54][71]=0;ram[54][72]=1;ram[54][73]=0;ram[54][74]=0;ram[54][75]=0;ram[54][76]=0;ram[54][77]=0;ram[54][78]=1;ram[54][79]=0;ram[54][80]=1;ram[54][81]=0;ram[54][82]=1;ram[54][83]=0;ram[54][84]=0;ram[54][85]=0;ram[54][86]=1;ram[54][87]=0;ram[54][88]=1;ram[54][89]=0;ram[54][90]=1;ram[54][91]=0;ram[54][92]=1;ram[54][93]=0;ram[54][94]=0;ram[54][95]=0;ram[54][96]=1;ram[54][97]=0;ram[54][98]=1;ram[54][99]=0;ram[54][100]=1;ram[54][101]=0;ram[54][102]=0;ram[54][103]=0;ram[54][104]=0;ram[54][105]=0;ram[54][106]=1;ram[54][107]=0;ram[54][108]=1;ram[54][109]=0;ram[54][110]=1;ram[54][111]=0;ram[54][112]=1;ram[54][113]=0;ram[54][114]=1;ram[54][115]=0;ram[54][116]=0;ram[54][117]=0;ram[54][118]=0;ram[54][119]=0;ram[54][120]=1;ram[54][121]=0;ram[54][122]=1;ram[54][123]=0;ram[54][124]=1;ram[54][125]=0;ram[54][126]=0;ram[54][127]=0;ram[54][128]=0;ram[54][129]=0;ram[54][130]=0;ram[54][131]=0;ram[54][132]=0;ram[54][133]=0;ram[54][134]=0;ram[54][135]=0;ram[54][136]=0;ram[54][137]=0;ram[54][138]=0;ram[54][139]=0;ram[54][140]=0;
        ram[55][0]=0;ram[55][1]=0;ram[55][2]=0;ram[55][3]=0;ram[55][4]=0;ram[55][5]=0;ram[55][6]=0;ram[55][7]=0;ram[55][8]=0;ram[55][9]=0;ram[55][10]=0;ram[55][11]=0;ram[55][12]=0;ram[55][13]=0;ram[55][14]=0;ram[55][15]=1;ram[55][16]=0;ram[55][17]=1;ram[55][18]=0;ram[55][19]=1;ram[55][20]=0;ram[55][21]=1;ram[55][22]=0;ram[55][23]=1;ram[55][24]=0;ram[55][25]=1;ram[55][26]=0;ram[55][27]=1;ram[55][28]=0;ram[55][29]=0;ram[55][30]=0;ram[55][31]=1;ram[55][32]=0;ram[55][33]=0;ram[55][34]=0;ram[55][35]=0;ram[55][36]=0;ram[55][37]=0;ram[55][38]=0;ram[55][39]=0;ram[55][40]=0;ram[55][41]=1;ram[55][42]=0;ram[55][43]=1;ram[55][44]=0;ram[55][45]=1;ram[55][46]=0;ram[55][47]=1;ram[55][48]=0;ram[55][49]=1;ram[55][50]=0;ram[55][51]=1;ram[55][52]=0;ram[55][53]=1;ram[55][54]=0;ram[55][55]=0;ram[55][56]=0;ram[55][57]=1;ram[55][58]=0;ram[55][59]=1;ram[55][60]=0;ram[55][61]=0;ram[55][62]=0;ram[55][63]=0;ram[55][64]=0;ram[55][65]=1;ram[55][66]=0;ram[55][67]=0;ram[55][68]=0;ram[55][69]=0;ram[55][70]=0;ram[55][71]=1;ram[55][72]=0;ram[55][73]=1;ram[55][74]=0;ram[55][75]=1;ram[55][76]=0;ram[55][77]=1;ram[55][78]=0;ram[55][79]=1;ram[55][80]=0;ram[55][81]=1;ram[55][82]=0;ram[55][83]=1;ram[55][84]=0;ram[55][85]=0;ram[55][86]=0;ram[55][87]=1;ram[55][88]=0;ram[55][89]=1;ram[55][90]=0;ram[55][91]=1;ram[55][92]=0;ram[55][93]=0;ram[55][94]=0;ram[55][95]=1;ram[55][96]=0;ram[55][97]=1;ram[55][98]=0;ram[55][99]=1;ram[55][100]=0;ram[55][101]=0;ram[55][102]=0;ram[55][103]=1;ram[55][104]=0;ram[55][105]=1;ram[55][106]=0;ram[55][107]=1;ram[55][108]=0;ram[55][109]=0;ram[55][110]=0;ram[55][111]=1;ram[55][112]=0;ram[55][113]=0;ram[55][114]=0;ram[55][115]=0;ram[55][116]=0;ram[55][117]=1;ram[55][118]=0;ram[55][119]=1;ram[55][120]=0;ram[55][121]=1;ram[55][122]=0;ram[55][123]=1;ram[55][124]=0;ram[55][125]=1;ram[55][126]=0;ram[55][127]=0;ram[55][128]=0;ram[55][129]=0;ram[55][130]=0;ram[55][131]=0;ram[55][132]=0;ram[55][133]=0;ram[55][134]=0;ram[55][135]=0;ram[55][136]=0;ram[55][137]=0;ram[55][138]=0;ram[55][139]=0;ram[55][140]=0;
        ram[56][0]=0;ram[56][1]=0;ram[56][2]=0;ram[56][3]=0;ram[56][4]=0;ram[56][5]=0;ram[56][6]=0;ram[56][7]=0;ram[56][8]=0;ram[56][9]=0;ram[56][10]=0;ram[56][11]=0;ram[56][12]=0;ram[56][13]=0;ram[56][14]=1;ram[56][15]=0;ram[56][16]=0;ram[56][17]=0;ram[56][18]=1;ram[56][19]=0;ram[56][20]=1;ram[56][21]=0;ram[56][22]=1;ram[56][23]=0;ram[56][24]=1;ram[56][25]=0;ram[56][26]=1;ram[56][27]=0;ram[56][28]=0;ram[56][29]=0;ram[56][30]=1;ram[56][31]=0;ram[56][32]=1;ram[56][33]=0;ram[56][34]=1;ram[56][35]=0;ram[56][36]=1;ram[56][37]=0;ram[56][38]=1;ram[56][39]=0;ram[56][40]=1;ram[56][41]=0;ram[56][42]=0;ram[56][43]=0;ram[56][44]=1;ram[56][45]=0;ram[56][46]=0;ram[56][47]=0;ram[56][48]=0;ram[56][49]=0;ram[56][50]=1;ram[56][51]=0;ram[56][52]=1;ram[56][53]=0;ram[56][54]=1;ram[56][55]=0;ram[56][56]=0;ram[56][57]=0;ram[56][58]=1;ram[56][59]=0;ram[56][60]=1;ram[56][61]=0;ram[56][62]=0;ram[56][63]=0;ram[56][64]=1;ram[56][65]=0;ram[56][66]=1;ram[56][67]=0;ram[56][68]=1;ram[56][69]=0;ram[56][70]=1;ram[56][71]=0;ram[56][72]=1;ram[56][73]=0;ram[56][74]=0;ram[56][75]=0;ram[56][76]=1;ram[56][77]=0;ram[56][78]=1;ram[56][79]=0;ram[56][80]=1;ram[56][81]=0;ram[56][82]=0;ram[56][83]=0;ram[56][84]=0;ram[56][85]=0;ram[56][86]=1;ram[56][87]=0;ram[56][88]=0;ram[56][89]=0;ram[56][90]=0;ram[56][91]=0;ram[56][92]=1;ram[56][93]=0;ram[56][94]=0;ram[56][95]=0;ram[56][96]=0;ram[56][97]=0;ram[56][98]=1;ram[56][99]=0;ram[56][100]=1;ram[56][101]=0;ram[56][102]=0;ram[56][103]=0;ram[56][104]=0;ram[56][105]=0;ram[56][106]=0;ram[56][107]=0;ram[56][108]=1;ram[56][109]=0;ram[56][110]=1;ram[56][111]=0;ram[56][112]=0;ram[56][113]=0;ram[56][114]=0;ram[56][115]=0;ram[56][116]=1;ram[56][117]=0;ram[56][118]=1;ram[56][119]=0;ram[56][120]=1;ram[56][121]=0;ram[56][122]=0;ram[56][123]=0;ram[56][124]=0;ram[56][125]=0;ram[56][126]=1;ram[56][127]=0;ram[56][128]=0;ram[56][129]=0;ram[56][130]=0;ram[56][131]=0;ram[56][132]=0;ram[56][133]=0;ram[56][134]=0;ram[56][135]=0;ram[56][136]=0;ram[56][137]=0;ram[56][138]=0;ram[56][139]=0;ram[56][140]=0;
        ram[57][0]=0;ram[57][1]=0;ram[57][2]=0;ram[57][3]=0;ram[57][4]=0;ram[57][5]=0;ram[57][6]=0;ram[57][7]=0;ram[57][8]=0;ram[57][9]=0;ram[57][10]=0;ram[57][11]=0;ram[57][12]=0;ram[57][13]=1;ram[57][14]=0;ram[57][15]=1;ram[57][16]=0;ram[57][17]=0;ram[57][18]=0;ram[57][19]=1;ram[57][20]=0;ram[57][21]=1;ram[57][22]=0;ram[57][23]=1;ram[57][24]=0;ram[57][25]=1;ram[57][26]=0;ram[57][27]=0;ram[57][28]=0;ram[57][29]=1;ram[57][30]=0;ram[57][31]=1;ram[57][32]=0;ram[57][33]=1;ram[57][34]=0;ram[57][35]=1;ram[57][36]=0;ram[57][37]=1;ram[57][38]=0;ram[57][39]=0;ram[57][40]=0;ram[57][41]=1;ram[57][42]=0;ram[57][43]=1;ram[57][44]=0;ram[57][45]=1;ram[57][46]=0;ram[57][47]=1;ram[57][48]=0;ram[57][49]=1;ram[57][50]=0;ram[57][51]=1;ram[57][52]=0;ram[57][53]=1;ram[57][54]=0;ram[57][55]=0;ram[57][56]=0;ram[57][57]=1;ram[57][58]=0;ram[57][59]=1;ram[57][60]=0;ram[57][61]=1;ram[57][62]=0;ram[57][63]=1;ram[57][64]=0;ram[57][65]=1;ram[57][66]=0;ram[57][67]=1;ram[57][68]=0;ram[57][69]=1;ram[57][70]=0;ram[57][71]=0;ram[57][72]=0;ram[57][73]=1;ram[57][74]=0;ram[57][75]=1;ram[57][76]=0;ram[57][77]=1;ram[57][78]=0;ram[57][79]=0;ram[57][80]=0;ram[57][81]=1;ram[57][82]=0;ram[57][83]=1;ram[57][84]=0;ram[57][85]=1;ram[57][86]=0;ram[57][87]=1;ram[57][88]=0;ram[57][89]=1;ram[57][90]=0;ram[57][91]=1;ram[57][92]=0;ram[57][93]=1;ram[57][94]=0;ram[57][95]=0;ram[57][96]=0;ram[57][97]=0;ram[57][98]=0;ram[57][99]=0;ram[57][100]=0;ram[57][101]=0;ram[57][102]=0;ram[57][103]=1;ram[57][104]=0;ram[57][105]=1;ram[57][106]=0;ram[57][107]=0;ram[57][108]=0;ram[57][109]=0;ram[57][110]=0;ram[57][111]=1;ram[57][112]=0;ram[57][113]=1;ram[57][114]=0;ram[57][115]=0;ram[57][116]=0;ram[57][117]=0;ram[57][118]=0;ram[57][119]=1;ram[57][120]=0;ram[57][121]=1;ram[57][122]=0;ram[57][123]=1;ram[57][124]=0;ram[57][125]=0;ram[57][126]=0;ram[57][127]=1;ram[57][128]=0;ram[57][129]=0;ram[57][130]=0;ram[57][131]=0;ram[57][132]=0;ram[57][133]=0;ram[57][134]=0;ram[57][135]=0;ram[57][136]=0;ram[57][137]=0;ram[57][138]=0;ram[57][139]=0;ram[57][140]=0;
        ram[58][0]=0;ram[58][1]=0;ram[58][2]=0;ram[58][3]=0;ram[58][4]=0;ram[58][5]=0;ram[58][6]=0;ram[58][7]=0;ram[58][8]=0;ram[58][9]=0;ram[58][10]=0;ram[58][11]=0;ram[58][12]=1;ram[58][13]=0;ram[58][14]=0;ram[58][15]=0;ram[58][16]=1;ram[58][17]=0;ram[58][18]=1;ram[58][19]=0;ram[58][20]=1;ram[58][21]=0;ram[58][22]=1;ram[58][23]=0;ram[58][24]=0;ram[58][25]=0;ram[58][26]=1;ram[58][27]=0;ram[58][28]=0;ram[58][29]=0;ram[58][30]=0;ram[58][31]=0;ram[58][32]=0;ram[58][33]=0;ram[58][34]=1;ram[58][35]=0;ram[58][36]=1;ram[58][37]=0;ram[58][38]=0;ram[58][39]=0;ram[58][40]=1;ram[58][41]=0;ram[58][42]=1;ram[58][43]=0;ram[58][44]=1;ram[58][45]=0;ram[58][46]=1;ram[58][47]=0;ram[58][48]=0;ram[58][49]=0;ram[58][50]=1;ram[58][51]=0;ram[58][52]=1;ram[58][53]=0;ram[58][54]=0;ram[58][55]=0;ram[58][56]=0;ram[58][57]=0;ram[58][58]=1;ram[58][59]=0;ram[58][60]=1;ram[58][61]=0;ram[58][62]=1;ram[58][63]=0;ram[58][64]=1;ram[58][65]=0;ram[58][66]=0;ram[58][67]=0;ram[58][68]=0;ram[58][69]=0;ram[58][70]=1;ram[58][71]=0;ram[58][72]=1;ram[58][73]=0;ram[58][74]=1;ram[58][75]=0;ram[58][76]=0;ram[58][77]=0;ram[58][78]=0;ram[58][79]=0;ram[58][80]=1;ram[58][81]=0;ram[58][82]=1;ram[58][83]=0;ram[58][84]=1;ram[58][85]=0;ram[58][86]=1;ram[58][87]=0;ram[58][88]=0;ram[58][89]=0;ram[58][90]=1;ram[58][91]=0;ram[58][92]=1;ram[58][93]=0;ram[58][94]=1;ram[58][95]=0;ram[58][96]=0;ram[58][97]=0;ram[58][98]=0;ram[58][99]=0;ram[58][100]=1;ram[58][101]=0;ram[58][102]=0;ram[58][103]=0;ram[58][104]=0;ram[58][105]=0;ram[58][106]=1;ram[58][107]=0;ram[58][108]=1;ram[58][109]=0;ram[58][110]=0;ram[58][111]=0;ram[58][112]=1;ram[58][113]=0;ram[58][114]=1;ram[58][115]=0;ram[58][116]=1;ram[58][117]=0;ram[58][118]=1;ram[58][119]=0;ram[58][120]=1;ram[58][121]=0;ram[58][122]=0;ram[58][123]=0;ram[58][124]=1;ram[58][125]=0;ram[58][126]=0;ram[58][127]=0;ram[58][128]=1;ram[58][129]=0;ram[58][130]=0;ram[58][131]=0;ram[58][132]=0;ram[58][133]=0;ram[58][134]=0;ram[58][135]=0;ram[58][136]=0;ram[58][137]=0;ram[58][138]=0;ram[58][139]=0;ram[58][140]=0;
        ram[59][0]=0;ram[59][1]=0;ram[59][2]=0;ram[59][3]=0;ram[59][4]=0;ram[59][5]=0;ram[59][6]=0;ram[59][7]=0;ram[59][8]=0;ram[59][9]=0;ram[59][10]=0;ram[59][11]=1;ram[59][12]=0;ram[59][13]=1;ram[59][14]=0;ram[59][15]=0;ram[59][16]=0;ram[59][17]=1;ram[59][18]=0;ram[59][19]=0;ram[59][20]=0;ram[59][21]=1;ram[59][22]=0;ram[59][23]=1;ram[59][24]=0;ram[59][25]=1;ram[59][26]=0;ram[59][27]=0;ram[59][28]=0;ram[59][29]=1;ram[59][30]=0;ram[59][31]=1;ram[59][32]=0;ram[59][33]=1;ram[59][34]=0;ram[59][35]=0;ram[59][36]=0;ram[59][37]=0;ram[59][38]=0;ram[59][39]=0;ram[59][40]=0;ram[59][41]=1;ram[59][42]=0;ram[59][43]=1;ram[59][44]=0;ram[59][45]=1;ram[59][46]=0;ram[59][47]=0;ram[59][48]=0;ram[59][49]=0;ram[59][50]=0;ram[59][51]=0;ram[59][52]=0;ram[59][53]=1;ram[59][54]=0;ram[59][55]=1;ram[59][56]=0;ram[59][57]=1;ram[59][58]=0;ram[59][59]=1;ram[59][60]=0;ram[59][61]=1;ram[59][62]=0;ram[59][63]=1;ram[59][64]=0;ram[59][65]=0;ram[59][66]=0;ram[59][67]=1;ram[59][68]=0;ram[59][69]=1;ram[59][70]=0;ram[59][71]=1;ram[59][72]=0;ram[59][73]=1;ram[59][74]=0;ram[59][75]=1;ram[59][76]=0;ram[59][77]=1;ram[59][78]=0;ram[59][79]=1;ram[59][80]=0;ram[59][81]=1;ram[59][82]=0;ram[59][83]=1;ram[59][84]=0;ram[59][85]=1;ram[59][86]=0;ram[59][87]=0;ram[59][88]=0;ram[59][89]=1;ram[59][90]=0;ram[59][91]=0;ram[59][92]=0;ram[59][93]=1;ram[59][94]=0;ram[59][95]=0;ram[59][96]=0;ram[59][97]=0;ram[59][98]=0;ram[59][99]=0;ram[59][100]=0;ram[59][101]=1;ram[59][102]=0;ram[59][103]=1;ram[59][104]=0;ram[59][105]=0;ram[59][106]=0;ram[59][107]=1;ram[59][108]=0;ram[59][109]=0;ram[59][110]=0;ram[59][111]=1;ram[59][112]=0;ram[59][113]=1;ram[59][114]=0;ram[59][115]=0;ram[59][116]=0;ram[59][117]=1;ram[59][118]=0;ram[59][119]=1;ram[59][120]=0;ram[59][121]=1;ram[59][122]=0;ram[59][123]=1;ram[59][124]=0;ram[59][125]=1;ram[59][126]=0;ram[59][127]=1;ram[59][128]=0;ram[59][129]=1;ram[59][130]=0;ram[59][131]=0;ram[59][132]=0;ram[59][133]=0;ram[59][134]=0;ram[59][135]=0;ram[59][136]=0;ram[59][137]=0;ram[59][138]=0;ram[59][139]=0;ram[59][140]=0;
        ram[60][0]=0;ram[60][1]=0;ram[60][2]=0;ram[60][3]=0;ram[60][4]=0;ram[60][5]=0;ram[60][6]=0;ram[60][7]=0;ram[60][8]=0;ram[60][9]=0;ram[60][10]=1;ram[60][11]=0;ram[60][12]=0;ram[60][13]=0;ram[60][14]=1;ram[60][15]=0;ram[60][16]=0;ram[60][17]=0;ram[60][18]=1;ram[60][19]=0;ram[60][20]=0;ram[60][21]=0;ram[60][22]=1;ram[60][23]=0;ram[60][24]=1;ram[60][25]=0;ram[60][26]=1;ram[60][27]=0;ram[60][28]=1;ram[60][29]=0;ram[60][30]=0;ram[60][31]=0;ram[60][32]=1;ram[60][33]=0;ram[60][34]=0;ram[60][35]=0;ram[60][36]=0;ram[60][37]=0;ram[60][38]=1;ram[60][39]=0;ram[60][40]=1;ram[60][41]=0;ram[60][42]=0;ram[60][43]=0;ram[60][44]=1;ram[60][45]=0;ram[60][46]=0;ram[60][47]=0;ram[60][48]=0;ram[60][49]=0;ram[60][50]=1;ram[60][51]=0;ram[60][52]=1;ram[60][53]=0;ram[60][54]=1;ram[60][55]=0;ram[60][56]=1;ram[60][57]=0;ram[60][58]=0;ram[60][59]=0;ram[60][60]=1;ram[60][61]=0;ram[60][62]=1;ram[60][63]=0;ram[60][64]=0;ram[60][65]=0;ram[60][66]=1;ram[60][67]=0;ram[60][68]=1;ram[60][69]=0;ram[60][70]=0;ram[60][71]=0;ram[60][72]=1;ram[60][73]=0;ram[60][74]=1;ram[60][75]=0;ram[60][76]=1;ram[60][77]=0;ram[60][78]=1;ram[60][79]=0;ram[60][80]=0;ram[60][81]=0;ram[60][82]=1;ram[60][83]=0;ram[60][84]=1;ram[60][85]=0;ram[60][86]=1;ram[60][87]=0;ram[60][88]=0;ram[60][89]=0;ram[60][90]=0;ram[60][91]=0;ram[60][92]=0;ram[60][93]=0;ram[60][94]=1;ram[60][95]=0;ram[60][96]=0;ram[60][97]=0;ram[60][98]=1;ram[60][99]=0;ram[60][100]=1;ram[60][101]=0;ram[60][102]=0;ram[60][103]=0;ram[60][104]=0;ram[60][105]=0;ram[60][106]=1;ram[60][107]=0;ram[60][108]=0;ram[60][109]=0;ram[60][110]=1;ram[60][111]=0;ram[60][112]=1;ram[60][113]=0;ram[60][114]=1;ram[60][115]=0;ram[60][116]=1;ram[60][117]=0;ram[60][118]=0;ram[60][119]=0;ram[60][120]=1;ram[60][121]=0;ram[60][122]=1;ram[60][123]=0;ram[60][124]=1;ram[60][125]=0;ram[60][126]=1;ram[60][127]=0;ram[60][128]=1;ram[60][129]=0;ram[60][130]=1;ram[60][131]=0;ram[60][132]=0;ram[60][133]=0;ram[60][134]=0;ram[60][135]=0;ram[60][136]=0;ram[60][137]=0;ram[60][138]=0;ram[60][139]=0;ram[60][140]=0;
        ram[61][0]=0;ram[61][1]=0;ram[61][2]=0;ram[61][3]=0;ram[61][4]=0;ram[61][5]=0;ram[61][6]=0;ram[61][7]=0;ram[61][8]=0;ram[61][9]=1;ram[61][10]=0;ram[61][11]=1;ram[61][12]=0;ram[61][13]=1;ram[61][14]=0;ram[61][15]=0;ram[61][16]=0;ram[61][17]=1;ram[61][18]=0;ram[61][19]=1;ram[61][20]=0;ram[61][21]=1;ram[61][22]=0;ram[61][23]=1;ram[61][24]=0;ram[61][25]=0;ram[61][26]=0;ram[61][27]=1;ram[61][28]=0;ram[61][29]=0;ram[61][30]=0;ram[61][31]=1;ram[61][32]=0;ram[61][33]=1;ram[61][34]=0;ram[61][35]=0;ram[61][36]=0;ram[61][37]=1;ram[61][38]=0;ram[61][39]=1;ram[61][40]=0;ram[61][41]=1;ram[61][42]=0;ram[61][43]=1;ram[61][44]=0;ram[61][45]=1;ram[61][46]=0;ram[61][47]=0;ram[61][48]=0;ram[61][49]=1;ram[61][50]=0;ram[61][51]=0;ram[61][52]=0;ram[61][53]=1;ram[61][54]=0;ram[61][55]=1;ram[61][56]=0;ram[61][57]=1;ram[61][58]=0;ram[61][59]=0;ram[61][60]=0;ram[61][61]=1;ram[61][62]=0;ram[61][63]=0;ram[61][64]=0;ram[61][65]=1;ram[61][66]=0;ram[61][67]=1;ram[61][68]=0;ram[61][69]=1;ram[61][70]=0;ram[61][71]=1;ram[61][72]=0;ram[61][73]=1;ram[61][74]=0;ram[61][75]=0;ram[61][76]=0;ram[61][77]=0;ram[61][78]=0;ram[61][79]=1;ram[61][80]=0;ram[61][81]=1;ram[61][82]=0;ram[61][83]=1;ram[61][84]=0;ram[61][85]=1;ram[61][86]=0;ram[61][87]=1;ram[61][88]=0;ram[61][89]=1;ram[61][90]=0;ram[61][91]=1;ram[61][92]=0;ram[61][93]=1;ram[61][94]=0;ram[61][95]=0;ram[61][96]=0;ram[61][97]=0;ram[61][98]=0;ram[61][99]=1;ram[61][100]=0;ram[61][101]=1;ram[61][102]=0;ram[61][103]=1;ram[61][104]=0;ram[61][105]=1;ram[61][106]=0;ram[61][107]=0;ram[61][108]=0;ram[61][109]=1;ram[61][110]=0;ram[61][111]=1;ram[61][112]=0;ram[61][113]=1;ram[61][114]=0;ram[61][115]=1;ram[61][116]=0;ram[61][117]=1;ram[61][118]=0;ram[61][119]=1;ram[61][120]=0;ram[61][121]=1;ram[61][122]=0;ram[61][123]=0;ram[61][124]=0;ram[61][125]=1;ram[61][126]=0;ram[61][127]=1;ram[61][128]=0;ram[61][129]=1;ram[61][130]=0;ram[61][131]=1;ram[61][132]=0;ram[61][133]=0;ram[61][134]=0;ram[61][135]=0;ram[61][136]=0;ram[61][137]=0;ram[61][138]=0;ram[61][139]=0;ram[61][140]=0;
        ram[62][0]=0;ram[62][1]=0;ram[62][2]=0;ram[62][3]=0;ram[62][4]=0;ram[62][5]=0;ram[62][6]=0;ram[62][7]=0;ram[62][8]=1;ram[62][9]=0;ram[62][10]=1;ram[62][11]=0;ram[62][12]=1;ram[62][13]=0;ram[62][14]=1;ram[62][15]=0;ram[62][16]=0;ram[62][17]=0;ram[62][18]=1;ram[62][19]=0;ram[62][20]=0;ram[62][21]=0;ram[62][22]=0;ram[62][23]=0;ram[62][24]=1;ram[62][25]=0;ram[62][26]=1;ram[62][27]=0;ram[62][28]=1;ram[62][29]=0;ram[62][30]=1;ram[62][31]=0;ram[62][32]=1;ram[62][33]=0;ram[62][34]=1;ram[62][35]=0;ram[62][36]=1;ram[62][37]=0;ram[62][38]=1;ram[62][39]=0;ram[62][40]=1;ram[62][41]=0;ram[62][42]=1;ram[62][43]=0;ram[62][44]=1;ram[62][45]=0;ram[62][46]=0;ram[62][47]=0;ram[62][48]=1;ram[62][49]=0;ram[62][50]=1;ram[62][51]=0;ram[62][52]=1;ram[62][53]=0;ram[62][54]=1;ram[62][55]=0;ram[62][56]=1;ram[62][57]=0;ram[62][58]=1;ram[62][59]=0;ram[62][60]=1;ram[62][61]=0;ram[62][62]=0;ram[62][63]=0;ram[62][64]=1;ram[62][65]=0;ram[62][66]=1;ram[62][67]=0;ram[62][68]=1;ram[62][69]=0;ram[62][70]=1;ram[62][71]=0;ram[62][72]=0;ram[62][73]=0;ram[62][74]=1;ram[62][75]=0;ram[62][76]=1;ram[62][77]=0;ram[62][78]=1;ram[62][79]=0;ram[62][80]=1;ram[62][81]=0;ram[62][82]=0;ram[62][83]=0;ram[62][84]=1;ram[62][85]=0;ram[62][86]=1;ram[62][87]=0;ram[62][88]=0;ram[62][89]=0;ram[62][90]=0;ram[62][91]=0;ram[62][92]=1;ram[62][93]=0;ram[62][94]=0;ram[62][95]=0;ram[62][96]=1;ram[62][97]=0;ram[62][98]=0;ram[62][99]=0;ram[62][100]=1;ram[62][101]=0;ram[62][102]=1;ram[62][103]=0;ram[62][104]=1;ram[62][105]=0;ram[62][106]=0;ram[62][107]=0;ram[62][108]=1;ram[62][109]=0;ram[62][110]=0;ram[62][111]=0;ram[62][112]=1;ram[62][113]=0;ram[62][114]=0;ram[62][115]=0;ram[62][116]=0;ram[62][117]=0;ram[62][118]=1;ram[62][119]=0;ram[62][120]=1;ram[62][121]=0;ram[62][122]=1;ram[62][123]=0;ram[62][124]=1;ram[62][125]=0;ram[62][126]=1;ram[62][127]=0;ram[62][128]=1;ram[62][129]=0;ram[62][130]=1;ram[62][131]=0;ram[62][132]=1;ram[62][133]=0;ram[62][134]=0;ram[62][135]=0;ram[62][136]=0;ram[62][137]=0;ram[62][138]=0;ram[62][139]=0;ram[62][140]=0;
        ram[63][0]=0;ram[63][1]=0;ram[63][2]=0;ram[63][3]=0;ram[63][4]=0;ram[63][5]=0;ram[63][6]=0;ram[63][7]=1;ram[63][8]=0;ram[63][9]=1;ram[63][10]=0;ram[63][11]=0;ram[63][12]=0;ram[63][13]=0;ram[63][14]=0;ram[63][15]=1;ram[63][16]=0;ram[63][17]=1;ram[63][18]=0;ram[63][19]=1;ram[63][20]=0;ram[63][21]=1;ram[63][22]=0;ram[63][23]=0;ram[63][24]=0;ram[63][25]=1;ram[63][26]=0;ram[63][27]=1;ram[63][28]=0;ram[63][29]=0;ram[63][30]=0;ram[63][31]=0;ram[63][32]=0;ram[63][33]=0;ram[63][34]=0;ram[63][35]=1;ram[63][36]=0;ram[63][37]=0;ram[63][38]=0;ram[63][39]=0;ram[63][40]=0;ram[63][41]=0;ram[63][42]=0;ram[63][43]=0;ram[63][44]=0;ram[63][45]=1;ram[63][46]=0;ram[63][47]=1;ram[63][48]=0;ram[63][49]=1;ram[63][50]=0;ram[63][51]=1;ram[63][52]=0;ram[63][53]=1;ram[63][54]=0;ram[63][55]=1;ram[63][56]=0;ram[63][57]=1;ram[63][58]=0;ram[63][59]=1;ram[63][60]=0;ram[63][61]=1;ram[63][62]=0;ram[63][63]=0;ram[63][64]=0;ram[63][65]=1;ram[63][66]=0;ram[63][67]=0;ram[63][68]=0;ram[63][69]=1;ram[63][70]=0;ram[63][71]=1;ram[63][72]=0;ram[63][73]=1;ram[63][74]=0;ram[63][75]=1;ram[63][76]=0;ram[63][77]=1;ram[63][78]=0;ram[63][79]=1;ram[63][80]=0;ram[63][81]=0;ram[63][82]=0;ram[63][83]=1;ram[63][84]=0;ram[63][85]=1;ram[63][86]=0;ram[63][87]=1;ram[63][88]=0;ram[63][89]=1;ram[63][90]=0;ram[63][91]=1;ram[63][92]=0;ram[63][93]=0;ram[63][94]=0;ram[63][95]=1;ram[63][96]=0;ram[63][97]=1;ram[63][98]=0;ram[63][99]=0;ram[63][100]=0;ram[63][101]=1;ram[63][102]=0;ram[63][103]=0;ram[63][104]=0;ram[63][105]=1;ram[63][106]=0;ram[63][107]=1;ram[63][108]=0;ram[63][109]=1;ram[63][110]=0;ram[63][111]=1;ram[63][112]=0;ram[63][113]=1;ram[63][114]=0;ram[63][115]=1;ram[63][116]=0;ram[63][117]=0;ram[63][118]=0;ram[63][119]=0;ram[63][120]=0;ram[63][121]=1;ram[63][122]=0;ram[63][123]=1;ram[63][124]=0;ram[63][125]=1;ram[63][126]=0;ram[63][127]=1;ram[63][128]=0;ram[63][129]=1;ram[63][130]=0;ram[63][131]=1;ram[63][132]=0;ram[63][133]=1;ram[63][134]=0;ram[63][135]=0;ram[63][136]=0;ram[63][137]=0;ram[63][138]=0;ram[63][139]=0;ram[63][140]=0;
        ram[64][0]=0;ram[64][1]=0;ram[64][2]=0;ram[64][3]=0;ram[64][4]=0;ram[64][5]=0;ram[64][6]=1;ram[64][7]=0;ram[64][8]=0;ram[64][9]=0;ram[64][10]=1;ram[64][11]=0;ram[64][12]=1;ram[64][13]=0;ram[64][14]=1;ram[64][15]=0;ram[64][16]=1;ram[64][17]=0;ram[64][18]=1;ram[64][19]=0;ram[64][20]=0;ram[64][21]=0;ram[64][22]=1;ram[64][23]=0;ram[64][24]=1;ram[64][25]=0;ram[64][26]=1;ram[64][27]=0;ram[64][28]=0;ram[64][29]=0;ram[64][30]=0;ram[64][31]=0;ram[64][32]=1;ram[64][33]=0;ram[64][34]=1;ram[64][35]=0;ram[64][36]=0;ram[64][37]=0;ram[64][38]=0;ram[64][39]=0;ram[64][40]=0;ram[64][41]=0;ram[64][42]=0;ram[64][43]=0;ram[64][44]=1;ram[64][45]=0;ram[64][46]=0;ram[64][47]=0;ram[64][48]=0;ram[64][49]=0;ram[64][50]=1;ram[64][51]=0;ram[64][52]=1;ram[64][53]=0;ram[64][54]=1;ram[64][55]=0;ram[64][56]=0;ram[64][57]=0;ram[64][58]=1;ram[64][59]=0;ram[64][60]=0;ram[64][61]=0;ram[64][62]=1;ram[64][63]=0;ram[64][64]=1;ram[64][65]=0;ram[64][66]=1;ram[64][67]=0;ram[64][68]=0;ram[64][69]=0;ram[64][70]=1;ram[64][71]=0;ram[64][72]=1;ram[64][73]=0;ram[64][74]=1;ram[64][75]=0;ram[64][76]=1;ram[64][77]=0;ram[64][78]=0;ram[64][79]=0;ram[64][80]=1;ram[64][81]=0;ram[64][82]=0;ram[64][83]=0;ram[64][84]=0;ram[64][85]=0;ram[64][86]=1;ram[64][87]=0;ram[64][88]=1;ram[64][89]=0;ram[64][90]=1;ram[64][91]=0;ram[64][92]=1;ram[64][93]=0;ram[64][94]=1;ram[64][95]=0;ram[64][96]=1;ram[64][97]=0;ram[64][98]=1;ram[64][99]=0;ram[64][100]=0;ram[64][101]=0;ram[64][102]=0;ram[64][103]=0;ram[64][104]=0;ram[64][105]=0;ram[64][106]=1;ram[64][107]=0;ram[64][108]=0;ram[64][109]=0;ram[64][110]=1;ram[64][111]=0;ram[64][112]=0;ram[64][113]=0;ram[64][114]=0;ram[64][115]=0;ram[64][116]=1;ram[64][117]=0;ram[64][118]=1;ram[64][119]=0;ram[64][120]=1;ram[64][121]=0;ram[64][122]=1;ram[64][123]=0;ram[64][124]=1;ram[64][125]=0;ram[64][126]=0;ram[64][127]=0;ram[64][128]=0;ram[64][129]=0;ram[64][130]=1;ram[64][131]=0;ram[64][132]=1;ram[64][133]=0;ram[64][134]=1;ram[64][135]=0;ram[64][136]=0;ram[64][137]=0;ram[64][138]=0;ram[64][139]=0;ram[64][140]=0;
        ram[65][0]=0;ram[65][1]=0;ram[65][2]=0;ram[65][3]=0;ram[65][4]=0;ram[65][5]=1;ram[65][6]=0;ram[65][7]=0;ram[65][8]=0;ram[65][9]=1;ram[65][10]=0;ram[65][11]=1;ram[65][12]=0;ram[65][13]=0;ram[65][14]=0;ram[65][15]=1;ram[65][16]=0;ram[65][17]=1;ram[65][18]=0;ram[65][19]=0;ram[65][20]=0;ram[65][21]=0;ram[65][22]=0;ram[65][23]=1;ram[65][24]=0;ram[65][25]=1;ram[65][26]=0;ram[65][27]=1;ram[65][28]=0;ram[65][29]=1;ram[65][30]=0;ram[65][31]=1;ram[65][32]=0;ram[65][33]=0;ram[65][34]=0;ram[65][35]=0;ram[65][36]=0;ram[65][37]=1;ram[65][38]=0;ram[65][39]=1;ram[65][40]=0;ram[65][41]=1;ram[65][42]=0;ram[65][43]=1;ram[65][44]=0;ram[65][45]=1;ram[65][46]=0;ram[65][47]=1;ram[65][48]=0;ram[65][49]=1;ram[65][50]=0;ram[65][51]=1;ram[65][52]=0;ram[65][53]=0;ram[65][54]=0;ram[65][55]=0;ram[65][56]=0;ram[65][57]=0;ram[65][58]=0;ram[65][59]=1;ram[65][60]=0;ram[65][61]=1;ram[65][62]=0;ram[65][63]=0;ram[65][64]=0;ram[65][65]=1;ram[65][66]=0;ram[65][67]=1;ram[65][68]=0;ram[65][69]=1;ram[65][70]=0;ram[65][71]=1;ram[65][72]=0;ram[65][73]=1;ram[65][74]=0;ram[65][75]=0;ram[65][76]=0;ram[65][77]=0;ram[65][78]=0;ram[65][79]=1;ram[65][80]=0;ram[65][81]=1;ram[65][82]=0;ram[65][83]=1;ram[65][84]=0;ram[65][85]=0;ram[65][86]=0;ram[65][87]=1;ram[65][88]=0;ram[65][89]=0;ram[65][90]=0;ram[65][91]=1;ram[65][92]=0;ram[65][93]=1;ram[65][94]=0;ram[65][95]=1;ram[65][96]=0;ram[65][97]=1;ram[65][98]=0;ram[65][99]=0;ram[65][100]=0;ram[65][101]=1;ram[65][102]=0;ram[65][103]=0;ram[65][104]=0;ram[65][105]=1;ram[65][106]=0;ram[65][107]=1;ram[65][108]=0;ram[65][109]=1;ram[65][110]=0;ram[65][111]=0;ram[65][112]=0;ram[65][113]=1;ram[65][114]=0;ram[65][115]=0;ram[65][116]=0;ram[65][117]=0;ram[65][118]=0;ram[65][119]=0;ram[65][120]=0;ram[65][121]=1;ram[65][122]=0;ram[65][123]=1;ram[65][124]=0;ram[65][125]=1;ram[65][126]=0;ram[65][127]=0;ram[65][128]=0;ram[65][129]=1;ram[65][130]=0;ram[65][131]=1;ram[65][132]=0;ram[65][133]=1;ram[65][134]=0;ram[65][135]=1;ram[65][136]=0;ram[65][137]=0;ram[65][138]=0;ram[65][139]=0;ram[65][140]=0;
        ram[66][0]=0;ram[66][1]=0;ram[66][2]=0;ram[66][3]=0;ram[66][4]=1;ram[66][5]=0;ram[66][6]=1;ram[66][7]=0;ram[66][8]=1;ram[66][9]=0;ram[66][10]=1;ram[66][11]=0;ram[66][12]=1;ram[66][13]=0;ram[66][14]=1;ram[66][15]=0;ram[66][16]=0;ram[66][17]=0;ram[66][18]=0;ram[66][19]=0;ram[66][20]=1;ram[66][21]=0;ram[66][22]=1;ram[66][23]=0;ram[66][24]=0;ram[66][25]=0;ram[66][26]=1;ram[66][27]=0;ram[66][28]=0;ram[66][29]=0;ram[66][30]=1;ram[66][31]=0;ram[66][32]=1;ram[66][33]=0;ram[66][34]=1;ram[66][35]=0;ram[66][36]=1;ram[66][37]=0;ram[66][38]=0;ram[66][39]=0;ram[66][40]=1;ram[66][41]=0;ram[66][42]=0;ram[66][43]=0;ram[66][44]=1;ram[66][45]=0;ram[66][46]=1;ram[66][47]=0;ram[66][48]=0;ram[66][49]=0;ram[66][50]=1;ram[66][51]=0;ram[66][52]=0;ram[66][53]=0;ram[66][54]=1;ram[66][55]=0;ram[66][56]=0;ram[66][57]=0;ram[66][58]=0;ram[66][59]=0;ram[66][60]=1;ram[66][61]=0;ram[66][62]=1;ram[66][63]=0;ram[66][64]=1;ram[66][65]=0;ram[66][66]=1;ram[66][67]=0;ram[66][68]=1;ram[66][69]=0;ram[66][70]=1;ram[66][71]=0;ram[66][72]=0;ram[66][73]=0;ram[66][74]=0;ram[66][75]=0;ram[66][76]=1;ram[66][77]=0;ram[66][78]=0;ram[66][79]=0;ram[66][80]=0;ram[66][81]=0;ram[66][82]=0;ram[66][83]=0;ram[66][84]=1;ram[66][85]=0;ram[66][86]=1;ram[66][87]=0;ram[66][88]=1;ram[66][89]=0;ram[66][90]=1;ram[66][91]=0;ram[66][92]=1;ram[66][93]=0;ram[66][94]=1;ram[66][95]=0;ram[66][96]=1;ram[66][97]=0;ram[66][98]=1;ram[66][99]=0;ram[66][100]=0;ram[66][101]=0;ram[66][102]=1;ram[66][103]=0;ram[66][104]=1;ram[66][105]=0;ram[66][106]=0;ram[66][107]=0;ram[66][108]=0;ram[66][109]=0;ram[66][110]=0;ram[66][111]=0;ram[66][112]=1;ram[66][113]=0;ram[66][114]=0;ram[66][115]=0;ram[66][116]=1;ram[66][117]=0;ram[66][118]=0;ram[66][119]=0;ram[66][120]=1;ram[66][121]=0;ram[66][122]=1;ram[66][123]=0;ram[66][124]=1;ram[66][125]=0;ram[66][126]=1;ram[66][127]=0;ram[66][128]=0;ram[66][129]=0;ram[66][130]=1;ram[66][131]=0;ram[66][132]=1;ram[66][133]=0;ram[66][134]=1;ram[66][135]=0;ram[66][136]=1;ram[66][137]=0;ram[66][138]=0;ram[66][139]=0;ram[66][140]=0;
        ram[67][0]=0;ram[67][1]=0;ram[67][2]=0;ram[67][3]=1;ram[67][4]=0;ram[67][5]=1;ram[67][6]=0;ram[67][7]=1;ram[67][8]=0;ram[67][9]=0;ram[67][10]=0;ram[67][11]=1;ram[67][12]=0;ram[67][13]=1;ram[67][14]=0;ram[67][15]=1;ram[67][16]=0;ram[67][17]=1;ram[67][18]=0;ram[67][19]=1;ram[67][20]=0;ram[67][21]=0;ram[67][22]=0;ram[67][23]=1;ram[67][24]=0;ram[67][25]=1;ram[67][26]=0;ram[67][27]=1;ram[67][28]=0;ram[67][29]=0;ram[67][30]=0;ram[67][31]=1;ram[67][32]=0;ram[67][33]=1;ram[67][34]=0;ram[67][35]=0;ram[67][36]=0;ram[67][37]=0;ram[67][38]=0;ram[67][39]=0;ram[67][40]=0;ram[67][41]=1;ram[67][42]=0;ram[67][43]=1;ram[67][44]=0;ram[67][45]=1;ram[67][46]=0;ram[67][47]=1;ram[67][48]=0;ram[67][49]=0;ram[67][50]=0;ram[67][51]=1;ram[67][52]=0;ram[67][53]=1;ram[67][54]=0;ram[67][55]=1;ram[67][56]=0;ram[67][57]=1;ram[67][58]=0;ram[67][59]=1;ram[67][60]=0;ram[67][61]=1;ram[67][62]=0;ram[67][63]=1;ram[67][64]=0;ram[67][65]=1;ram[67][66]=0;ram[67][67]=1;ram[67][68]=0;ram[67][69]=1;ram[67][70]=0;ram[67][71]=0;ram[67][72]=0;ram[67][73]=0;ram[67][74]=0;ram[67][75]=0;ram[67][76]=0;ram[67][77]=1;ram[67][78]=0;ram[67][79]=1;ram[67][80]=0;ram[67][81]=1;ram[67][82]=0;ram[67][83]=1;ram[67][84]=0;ram[67][85]=1;ram[67][86]=0;ram[67][87]=1;ram[67][88]=0;ram[67][89]=1;ram[67][90]=0;ram[67][91]=0;ram[67][92]=0;ram[67][93]=0;ram[67][94]=0;ram[67][95]=1;ram[67][96]=0;ram[67][97]=0;ram[67][98]=0;ram[67][99]=0;ram[67][100]=0;ram[67][101]=0;ram[67][102]=0;ram[67][103]=0;ram[67][104]=0;ram[67][105]=1;ram[67][106]=0;ram[67][107]=0;ram[67][108]=0;ram[67][109]=0;ram[67][110]=0;ram[67][111]=0;ram[67][112]=0;ram[67][113]=1;ram[67][114]=0;ram[67][115]=1;ram[67][116]=0;ram[67][117]=0;ram[67][118]=0;ram[67][119]=1;ram[67][120]=0;ram[67][121]=1;ram[67][122]=0;ram[67][123]=1;ram[67][124]=0;ram[67][125]=1;ram[67][126]=0;ram[67][127]=1;ram[67][128]=0;ram[67][129]=1;ram[67][130]=0;ram[67][131]=1;ram[67][132]=0;ram[67][133]=1;ram[67][134]=0;ram[67][135]=1;ram[67][136]=0;ram[67][137]=1;ram[67][138]=0;ram[67][139]=0;ram[67][140]=0;
        ram[68][0]=0;ram[68][1]=0;ram[68][2]=1;ram[68][3]=0;ram[68][4]=1;ram[68][5]=0;ram[68][6]=1;ram[68][7]=0;ram[68][8]=0;ram[68][9]=0;ram[68][10]=1;ram[68][11]=0;ram[68][12]=1;ram[68][13]=0;ram[68][14]=1;ram[68][15]=0;ram[68][16]=1;ram[68][17]=0;ram[68][18]=0;ram[68][19]=0;ram[68][20]=1;ram[68][21]=0;ram[68][22]=0;ram[68][23]=0;ram[68][24]=1;ram[68][25]=0;ram[68][26]=1;ram[68][27]=0;ram[68][28]=0;ram[68][29]=0;ram[68][30]=1;ram[68][31]=0;ram[68][32]=0;ram[68][33]=0;ram[68][34]=1;ram[68][35]=0;ram[68][36]=0;ram[68][37]=0;ram[68][38]=1;ram[68][39]=0;ram[68][40]=1;ram[68][41]=0;ram[68][42]=1;ram[68][43]=0;ram[68][44]=1;ram[68][45]=0;ram[68][46]=0;ram[68][47]=0;ram[68][48]=0;ram[68][49]=0;ram[68][50]=1;ram[68][51]=0;ram[68][52]=1;ram[68][53]=0;ram[68][54]=0;ram[68][55]=0;ram[68][56]=1;ram[68][57]=0;ram[68][58]=0;ram[68][59]=0;ram[68][60]=0;ram[68][61]=0;ram[68][62]=1;ram[68][63]=0;ram[68][64]=0;ram[68][65]=0;ram[68][66]=1;ram[68][67]=0;ram[68][68]=1;ram[68][69]=0;ram[68][70]=0;ram[68][71]=0;ram[68][72]=1;ram[68][73]=0;ram[68][74]=1;ram[68][75]=0;ram[68][76]=1;ram[68][77]=0;ram[68][78]=1;ram[68][79]=0;ram[68][80]=1;ram[68][81]=0;ram[68][82]=0;ram[68][83]=0;ram[68][84]=1;ram[68][85]=0;ram[68][86]=0;ram[68][87]=0;ram[68][88]=1;ram[68][89]=0;ram[68][90]=0;ram[68][91]=0;ram[68][92]=1;ram[68][93]=0;ram[68][94]=1;ram[68][95]=0;ram[68][96]=1;ram[68][97]=0;ram[68][98]=1;ram[68][99]=0;ram[68][100]=1;ram[68][101]=0;ram[68][102]=1;ram[68][103]=0;ram[68][104]=0;ram[68][105]=0;ram[68][106]=1;ram[68][107]=0;ram[68][108]=0;ram[68][109]=0;ram[68][110]=1;ram[68][111]=0;ram[68][112]=1;ram[68][113]=0;ram[68][114]=1;ram[68][115]=0;ram[68][116]=0;ram[68][117]=0;ram[68][118]=0;ram[68][119]=0;ram[68][120]=1;ram[68][121]=0;ram[68][122]=1;ram[68][123]=0;ram[68][124]=1;ram[68][125]=0;ram[68][126]=1;ram[68][127]=0;ram[68][128]=0;ram[68][129]=0;ram[68][130]=0;ram[68][131]=0;ram[68][132]=1;ram[68][133]=0;ram[68][134]=1;ram[68][135]=0;ram[68][136]=1;ram[68][137]=0;ram[68][138]=1;ram[68][139]=0;ram[68][140]=0;
        ram[69][0]=0;ram[69][1]=1;ram[69][2]=0;ram[69][3]=0;ram[69][4]=0;ram[69][5]=0;ram[69][6]=0;ram[69][7]=1;ram[69][8]=0;ram[69][9]=1;ram[69][10]=0;ram[69][11]=1;ram[69][12]=0;ram[69][13]=1;ram[69][14]=0;ram[69][15]=1;ram[69][16]=0;ram[69][17]=1;ram[69][18]=0;ram[69][19]=0;ram[69][20]=0;ram[69][21]=0;ram[69][22]=0;ram[69][23]=0;ram[69][24]=0;ram[69][25]=1;ram[69][26]=0;ram[69][27]=1;ram[69][28]=0;ram[69][29]=0;ram[69][30]=0;ram[69][31]=0;ram[69][32]=0;ram[69][33]=1;ram[69][34]=0;ram[69][35]=1;ram[69][36]=0;ram[69][37]=1;ram[69][38]=0;ram[69][39]=1;ram[69][40]=0;ram[69][41]=1;ram[69][42]=0;ram[69][43]=1;ram[69][44]=0;ram[69][45]=0;ram[69][46]=0;ram[69][47]=1;ram[69][48]=0;ram[69][49]=0;ram[69][50]=0;ram[69][51]=0;ram[69][52]=0;ram[69][53]=0;ram[69][54]=0;ram[69][55]=1;ram[69][56]=0;ram[69][57]=1;ram[69][58]=0;ram[69][59]=0;ram[69][60]=0;ram[69][61]=0;ram[69][62]=0;ram[69][63]=1;ram[69][64]=0;ram[69][65]=1;ram[69][66]=0;ram[69][67]=1;ram[69][68]=0;ram[69][69]=0;ram[69][70]=0;ram[69][71]=1;ram[69][72]=0;ram[69][73]=1;ram[69][74]=0;ram[69][75]=0;ram[69][76]=0;ram[69][77]=1;ram[69][78]=0;ram[69][79]=1;ram[69][80]=0;ram[69][81]=0;ram[69][82]=0;ram[69][83]=0;ram[69][84]=0;ram[69][85]=1;ram[69][86]=0;ram[69][87]=1;ram[69][88]=0;ram[69][89]=0;ram[69][90]=0;ram[69][91]=1;ram[69][92]=0;ram[69][93]=1;ram[69][94]=0;ram[69][95]=0;ram[69][96]=0;ram[69][97]=1;ram[69][98]=0;ram[69][99]=1;ram[69][100]=0;ram[69][101]=0;ram[69][102]=0;ram[69][103]=0;ram[69][104]=0;ram[69][105]=0;ram[69][106]=0;ram[69][107]=0;ram[69][108]=0;ram[69][109]=0;ram[69][110]=0;ram[69][111]=1;ram[69][112]=0;ram[69][113]=1;ram[69][114]=0;ram[69][115]=1;ram[69][116]=0;ram[69][117]=1;ram[69][118]=0;ram[69][119]=0;ram[69][120]=0;ram[69][121]=1;ram[69][122]=0;ram[69][123]=1;ram[69][124]=0;ram[69][125]=0;ram[69][126]=0;ram[69][127]=0;ram[69][128]=0;ram[69][129]=1;ram[69][130]=0;ram[69][131]=0;ram[69][132]=0;ram[69][133]=1;ram[69][134]=0;ram[69][135]=0;ram[69][136]=0;ram[69][137]=0;ram[69][138]=0;ram[69][139]=1;ram[69][140]=0;
        
        ans2_ram[0]<=0;ans2_ram[1]<=0;ans2_ram[2]<=0;ans2_ram[3]<=0;ans2_ram[4]<=0;ans2_ram[5]<=0;ans2_ram[6]<=0;ans2_ram[7]<=0;ans2_ram[8]<=0;ans2_ram[9]<=0;ans2_ram[10]<=0;ans2_ram[11]<=0;ans2_ram[12]<=0;ans2_ram[13]<=0;ans2_ram[14]<=0;ans2_ram[15]<=0;ans2_ram[16]<=0;ans2_ram[17]<=0;ans2_ram[18]<=0;ans2_ram[19]<=0;ans2_ram[20]<=0;ans2_ram[21]<=0;ans2_ram[22]<=0;ans2_ram[23]<=0;ans2_ram[24]<=0;ans2_ram[25]<=0;ans2_ram[26]<=0;ans2_ram[27]<=0;ans2_ram[28]<=0;ans2_ram[29]<=0;ans2_ram[30]<=0;ans2_ram[31]<=0;ans2_ram[32]<=0;ans2_ram[33]<=0;ans2_ram[34]<=0;ans2_ram[35]<=0;ans2_ram[36]<=0;ans2_ram[37]<=0;ans2_ram[38]<=0;ans2_ram[39]<=0;ans2_ram[40]<=0;ans2_ram[41]<=0;ans2_ram[42]<=0;ans2_ram[43]<=0;ans2_ram[44]<=0;ans2_ram[45]<=0;ans2_ram[46]<=0;ans2_ram[47]<=0;ans2_ram[48]<=0;ans2_ram[49]<=0;ans2_ram[50]<=0;ans2_ram[51]<=0;ans2_ram[52]<=0;ans2_ram[53]<=0;ans2_ram[54]<=0;ans2_ram[55]<=0;ans2_ram[56]<=0;ans2_ram[57]<=0;ans2_ram[58]<=0;ans2_ram[59]<=0;ans2_ram[60]<=0;ans2_ram[61]<=0;ans2_ram[62]<=0;ans2_ram[63]<=0;ans2_ram[64]<=0;ans2_ram[65]<=0;ans2_ram[66]<=0;ans2_ram[67]<=0;ans2_ram[68]<=0;ans2_ram[69]<=0;
        ans2_ram[70]<=1;
        ans2_ram[71]<=0;ans2_ram[72]<=0;ans2_ram[73]<=0;ans2_ram[74]<=0;ans2_ram[75]<=0;ans2_ram[76]<=0;ans2_ram[77]<=0;ans2_ram[78]<=0;ans2_ram[79]<=0;ans2_ram[80]<=0;ans2_ram[81]<=0;ans2_ram[82]<=0;ans2_ram[83]<=0;ans2_ram[84]<=0;ans2_ram[85]<=0;ans2_ram[86]<=0;ans2_ram[87]<=0;ans2_ram[88]<=0;ans2_ram[89]<=0;ans2_ram[90]<=0;ans2_ram[91]<=0;ans2_ram[92]<=0;ans2_ram[93]<=0;ans2_ram[94]<=0;ans2_ram[95]<=0;ans2_ram[96]<=0;ans2_ram[97]<=0;ans2_ram[98]<=0;ans2_ram[99]<=0;ans2_ram[100]<=0;ans2_ram[101]<=0;ans2_ram[102]<=0;ans2_ram[103]<=0;ans2_ram[104]<=0;ans2_ram[105]<=0;ans2_ram[106]<=0;ans2_ram[107]<=0;ans2_ram[108]<=0;ans2_ram[109]<=0;ans2_ram[110]<=0;ans2_ram[111]<=0;ans2_ram[112]<=0;ans2_ram[113]<=0;ans2_ram[114]<=0;ans2_ram[115]<=0;ans2_ram[116]<=0;ans2_ram[117]<=0;ans2_ram[118]<=0;ans2_ram[119]<=0;ans2_ram[120]<=0;ans2_ram[121]<=0;ans2_ram[122]<=0;ans2_ram[123]<=0;ans2_ram[124]<=0;ans2_ram[125]<=0;ans2_ram[126]<=0;ans2_ram[127]<=0;ans2_ram[128]<=0;ans2_ram[129]<=0;ans2_ram[130]<=0;ans2_ram[131]<=0;ans2_ram[132]<=0;ans2_ram[133]<=0;ans2_ram[134]<=0;ans2_ram[135]<=0;ans2_ram[136]<=0;ans2_ram[137]<=0;ans2_ram[138]<=0;ans2_ram[139]<=0;ans2_ram[140]<=0;
        
        ans1=0;ans2=0;
    end
    
    reg [7:0]pos=0;
    always @(posedge clk)
    begin
        if(rst)pos<=0;
        else if (pos<size/2-1)pos<=pos+1;
    end
    
    reg [size-1:0]compare={{70{1'b0}},1'b1,{70{1'b0}}};
    genvar i;
    generate
        for(i=0;i<size;i=i+1)
        begin: To_The_Moon
            if(i==0)
            begin
                always @(posedge clk)
                begin
                    if (rst || ram[pos][i])
                    begin
                        compare[i]<=0;
                        ans2_ram[i]<=0;
                    end
                    else if (ram[pos][i+1] && compare[i+1])
                    begin
                        compare[i]<=1;
                        ans2_ram[i]<=ans2_ram[i]+ans2_ram[i+1];
                    end
                end
            end
            else if(i==size-1)
            begin
                always @(posedge clk)
                begin
                    if (rst || ram[pos][i])
                    begin
                        compare[i]<=0;
                        ans2_ram[i]<=0;
                    end
                    else if (ram[pos][i-1] && compare[i-1])
                    begin
                        compare[i]<=1;
                        ans2_ram[i]<=ans2_ram[i]+ans2_ram[i-1];
                    end
                end
            end
            else
            begin
                always @(posedge clk)
                begin
                    if (rst || ram[pos][i])
                    begin
                        compare[i]<=0;
                        ans2_ram[i]<=0;
                    end
                    else if ((ram[pos][i+1] && compare[i+1]) && (ram[pos][i-1] && compare[i-1]))
                    begin
                        compare[i]<=1;
                        ans2_ram[i]<=ans2_ram[i]+ans2_ram[i-1]+ans2_ram[i+1];
                    end
                    else if (ram[pos][i+1] && compare[i+1])
                    begin
                        compare[i]<=1;
                        ans2_ram[i]<=ans2_ram[i]+ans2_ram[i+1];
                    end
                    else if (ram[pos][i-1] && compare[i-1])
                    begin
                        compare[i]<=1;
                        ans2_ram[i]<=ans2_ram[i]+ans2_ram[i-1];
                    end
                end
            end
        end
    endgenerate
    
    integer j=0;
    always @(posedge clk)
    begin
        if(rst || pos>size/2-1) 
        begin
            ans1<=0;
        end
        else
        begin
            for(j=0;j<size;j=j+1) 
            begin
                ans1=ans1+(ram[pos][j]&&compare[j]);
            end
        end
    end
    
    integer k=0;
    always @(*)
    begin
        ans2=0;
        for (k=0;k<size;k=k+1)
        begin: add_ans2
            ans2=ans2+ans2_ram[k];
        end
    end
    
endmodule
