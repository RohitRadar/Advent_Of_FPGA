`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.01.2026 10:08:04
// Design Name: 
// Module Name: Main2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Main2(
    input clk,rst,
    output reg [31:0]sum
    );
    parameter size=137;
    
    reg [size-1:0]ram[size-1:0];
    reg [size-1:0]sumram[size-1:0];
    initial
    begin
        ram[0][0]=1;ram[0][1]=1;ram[0][2]=0;ram[0][3]=1;ram[0][4]=1;ram[0][5]=1;ram[0][6]=1;ram[0][7]=0;ram[0][8]=0;ram[0][9]=1;ram[0][10]=1;ram[0][11]=1;ram[0][12]=0;ram[0][13]=0;ram[0][14]=1;ram[0][15]=1;ram[0][16]=1;ram[0][17]=0;ram[0][18]=1;ram[0][19]=1;ram[0][20]=0;ram[0][21]=1;ram[0][22]=1;ram[0][23]=1;ram[0][24]=1;ram[0][25]=1;ram[0][26]=1;ram[0][27]=1;ram[0][28]=0;ram[0][29]=1;ram[0][30]=1;ram[0][31]=1;ram[0][32]=0;ram[0][33]=1;ram[0][34]=1;ram[0][35]=1;ram[0][36]=1;ram[0][37]=1;ram[0][38]=1;ram[0][39]=1;ram[0][40]=1;ram[0][41]=0;ram[0][42]=1;ram[0][43]=1;ram[0][44]=1;ram[0][45]=1;ram[0][46]=1;ram[0][47]=1;ram[0][48]=1;ram[0][49]=0;ram[0][50]=0;ram[0][51]=1;ram[0][52]=1;ram[0][53]=1;ram[0][54]=1;ram[0][55]=1;ram[0][56]=1;ram[0][57]=0;ram[0][58]=1;ram[0][59]=1;ram[0][60]=0;ram[0][61]=0;ram[0][62]=0;ram[0][63]=0;ram[0][64]=0;ram[0][65]=1;ram[0][66]=1;ram[0][67]=0;ram[0][68]=1;ram[0][69]=0;ram[0][70]=0;ram[0][71]=1;ram[0][72]=0;ram[0][73]=1;ram[0][74]=1;ram[0][75]=1;ram[0][76]=0;ram[0][77]=1;ram[0][78]=0;ram[0][79]=1;ram[0][80]=0;ram[0][81]=1;ram[0][82]=1;ram[0][83]=1;ram[0][84]=0;ram[0][85]=1;ram[0][86]=0;ram[0][87]=0;ram[0][88]=0;ram[0][89]=1;ram[0][90]=1;ram[0][91]=1;ram[0][92]=1;ram[0][93]=1;ram[0][94]=0;ram[0][95]=1;ram[0][96]=0;ram[0][97]=1;ram[0][98]=0;ram[0][99]=1;ram[0][100]=0;ram[0][101]=1;ram[0][102]=0;ram[0][103]=1;ram[0][104]=1;ram[0][105]=1;ram[0][106]=1;ram[0][107]=1;ram[0][108]=1;ram[0][109]=1;ram[0][110]=0;ram[0][111]=0;ram[0][112]=0;ram[0][113]=1;ram[0][114]=0;ram[0][115]=0;ram[0][116]=0;ram[0][117]=1;ram[0][118]=0;ram[0][119]=1;ram[0][120]=0;ram[0][121]=0;ram[0][122]=0;ram[0][123]=1;ram[0][124]=0;ram[0][125]=1;ram[0][126]=0;ram[0][127]=1;ram[0][128]=1;ram[0][129]=1;ram[0][130]=1;ram[0][131]=1;ram[0][132]=1;ram[0][133]=1;ram[0][134]=1;ram[0][135]=1;ram[0][136]=1;
        ram[1][0]=0;ram[1][1]=1;ram[1][2]=0;ram[1][3]=1;ram[1][4]=1;ram[1][5]=0;ram[1][6]=1;ram[1][7]=1;ram[1][8]=0;ram[1][9]=0;ram[1][10]=1;ram[1][11]=1;ram[1][12]=1;ram[1][13]=1;ram[1][14]=1;ram[1][15]=0;ram[1][16]=1;ram[1][17]=0;ram[1][18]=0;ram[1][19]=1;ram[1][20]=0;ram[1][21]=0;ram[1][22]=1;ram[1][23]=1;ram[1][24]=0;ram[1][25]=0;ram[1][26]=1;ram[1][27]=1;ram[1][28]=0;ram[1][29]=1;ram[1][30]=1;ram[1][31]=1;ram[1][32]=0;ram[1][33]=1;ram[1][34]=1;ram[1][35]=0;ram[1][36]=0;ram[1][37]=0;ram[1][38]=1;ram[1][39]=1;ram[1][40]=0;ram[1][41]=1;ram[1][42]=0;ram[1][43]=1;ram[1][44]=0;ram[1][45]=1;ram[1][46]=0;ram[1][47]=1;ram[1][48]=0;ram[1][49]=0;ram[1][50]=1;ram[1][51]=0;ram[1][52]=0;ram[1][53]=1;ram[1][54]=1;ram[1][55]=0;ram[1][56]=1;ram[1][57]=1;ram[1][58]=1;ram[1][59]=1;ram[1][60]=0;ram[1][61]=1;ram[1][62]=0;ram[1][63]=1;ram[1][64]=1;ram[1][65]=1;ram[1][66]=1;ram[1][67]=1;ram[1][68]=1;ram[1][69]=1;ram[1][70]=1;ram[1][71]=0;ram[1][72]=1;ram[1][73]=1;ram[1][74]=0;ram[1][75]=1;ram[1][76]=0;ram[1][77]=1;ram[1][78]=0;ram[1][79]=1;ram[1][80]=0;ram[1][81]=1;ram[1][82]=1;ram[1][83]=1;ram[1][84]=0;ram[1][85]=0;ram[1][86]=1;ram[1][87]=1;ram[1][88]=1;ram[1][89]=1;ram[1][90]=1;ram[1][91]=0;ram[1][92]=0;ram[1][93]=1;ram[1][94]=0;ram[1][95]=1;ram[1][96]=1;ram[1][97]=1;ram[1][98]=0;ram[1][99]=1;ram[1][100]=0;ram[1][101]=1;ram[1][102]=0;ram[1][103]=0;ram[1][104]=1;ram[1][105]=1;ram[1][106]=0;ram[1][107]=0;ram[1][108]=1;ram[1][109]=1;ram[1][110]=0;ram[1][111]=1;ram[1][112]=1;ram[1][113]=1;ram[1][114]=0;ram[1][115]=1;ram[1][116]=0;ram[1][117]=0;ram[1][118]=0;ram[1][119]=1;ram[1][120]=1;ram[1][121]=0;ram[1][122]=1;ram[1][123]=1;ram[1][124]=1;ram[1][125]=1;ram[1][126]=1;ram[1][127]=0;ram[1][128]=1;ram[1][129]=0;ram[1][130]=0;ram[1][131]=1;ram[1][132]=0;ram[1][133]=0;ram[1][134]=1;ram[1][135]=0;ram[1][136]=1;
        ram[2][0]=0;ram[2][1]=1;ram[2][2]=0;ram[2][3]=1;ram[2][4]=1;ram[2][5]=1;ram[2][6]=0;ram[2][7]=1;ram[2][8]=1;ram[2][9]=0;ram[2][10]=1;ram[2][11]=0;ram[2][12]=1;ram[2][13]=1;ram[2][14]=0;ram[2][15]=1;ram[2][16]=1;ram[2][17]=1;ram[2][18]=1;ram[2][19]=1;ram[2][20]=0;ram[2][21]=1;ram[2][22]=0;ram[2][23]=1;ram[2][24]=1;ram[2][25]=1;ram[2][26]=0;ram[2][27]=1;ram[2][28]=0;ram[2][29]=1;ram[2][30]=1;ram[2][31]=1;ram[2][32]=1;ram[2][33]=1;ram[2][34]=0;ram[2][35]=1;ram[2][36]=0;ram[2][37]=0;ram[2][38]=0;ram[2][39]=1;ram[2][40]=1;ram[2][41]=1;ram[2][42]=1;ram[2][43]=1;ram[2][44]=1;ram[2][45]=1;ram[2][46]=1;ram[2][47]=1;ram[2][48]=0;ram[2][49]=1;ram[2][50]=1;ram[2][51]=1;ram[2][52]=0;ram[2][53]=1;ram[2][54]=1;ram[2][55]=0;ram[2][56]=1;ram[2][57]=1;ram[2][58]=0;ram[2][59]=1;ram[2][60]=0;ram[2][61]=0;ram[2][62]=1;ram[2][63]=1;ram[2][64]=0;ram[2][65]=0;ram[2][66]=1;ram[2][67]=0;ram[2][68]=1;ram[2][69]=1;ram[2][70]=1;ram[2][71]=1;ram[2][72]=0;ram[2][73]=0;ram[2][74]=1;ram[2][75]=1;ram[2][76]=1;ram[2][77]=0;ram[2][78]=0;ram[2][79]=0;ram[2][80]=1;ram[2][81]=0;ram[2][82]=1;ram[2][83]=0;ram[2][84]=1;ram[2][85]=1;ram[2][86]=1;ram[2][87]=1;ram[2][88]=0;ram[2][89]=0;ram[2][90]=1;ram[2][91]=0;ram[2][92]=0;ram[2][93]=1;ram[2][94]=1;ram[2][95]=0;ram[2][96]=1;ram[2][97]=1;ram[2][98]=0;ram[2][99]=0;ram[2][100]=0;ram[2][101]=1;ram[2][102]=0;ram[2][103]=1;ram[2][104]=0;ram[2][105]=0;ram[2][106]=1;ram[2][107]=1;ram[2][108]=1;ram[2][109]=1;ram[2][110]=1;ram[2][111]=1;ram[2][112]=1;ram[2][113]=0;ram[2][114]=1;ram[2][115]=1;ram[2][116]=1;ram[2][117]=0;ram[2][118]=0;ram[2][119]=1;ram[2][120]=1;ram[2][121]=1;ram[2][122]=0;ram[2][123]=0;ram[2][124]=1;ram[2][125]=1;ram[2][126]=1;ram[2][127]=1;ram[2][128]=0;ram[2][129]=1;ram[2][130]=1;ram[2][131]=1;ram[2][132]=0;ram[2][133]=1;ram[2][134]=1;ram[2][135]=1;ram[2][136]=1;
        ram[3][0]=1;ram[3][1]=1;ram[3][2]=0;ram[3][3]=1;ram[3][4]=1;ram[3][5]=1;ram[3][6]=1;ram[3][7]=1;ram[3][8]=1;ram[3][9]=0;ram[3][10]=1;ram[3][11]=1;ram[3][12]=1;ram[3][13]=0;ram[3][14]=0;ram[3][15]=0;ram[3][16]=1;ram[3][17]=1;ram[3][18]=0;ram[3][19]=1;ram[3][20]=1;ram[3][21]=1;ram[3][22]=0;ram[3][23]=0;ram[3][24]=1;ram[3][25]=1;ram[3][26]=1;ram[3][27]=0;ram[3][28]=0;ram[3][29]=0;ram[3][30]=0;ram[3][31]=1;ram[3][32]=0;ram[3][33]=1;ram[3][34]=1;ram[3][35]=1;ram[3][36]=1;ram[3][37]=1;ram[3][38]=1;ram[3][39]=0;ram[3][40]=1;ram[3][41]=1;ram[3][42]=1;ram[3][43]=0;ram[3][44]=1;ram[3][45]=0;ram[3][46]=0;ram[3][47]=1;ram[3][48]=0;ram[3][49]=0;ram[3][50]=1;ram[3][51]=1;ram[3][52]=1;ram[3][53]=0;ram[3][54]=1;ram[3][55]=1;ram[3][56]=0;ram[3][57]=0;ram[3][58]=0;ram[3][59]=0;ram[3][60]=1;ram[3][61]=0;ram[3][62]=0;ram[3][63]=0;ram[3][64]=1;ram[3][65]=1;ram[3][66]=1;ram[3][67]=0;ram[3][68]=1;ram[3][69]=1;ram[3][70]=0;ram[3][71]=0;ram[3][72]=1;ram[3][73]=0;ram[3][74]=1;ram[3][75]=1;ram[3][76]=1;ram[3][77]=1;ram[3][78]=0;ram[3][79]=0;ram[3][80]=1;ram[3][81]=1;ram[3][82]=1;ram[3][83]=0;ram[3][84]=0;ram[3][85]=0;ram[3][86]=1;ram[3][87]=1;ram[3][88]=0;ram[3][89]=1;ram[3][90]=0;ram[3][91]=0;ram[3][92]=1;ram[3][93]=1;ram[3][94]=0;ram[3][95]=1;ram[3][96]=1;ram[3][97]=1;ram[3][98]=0;ram[3][99]=0;ram[3][100]=0;ram[3][101]=1;ram[3][102]=0;ram[3][103]=1;ram[3][104]=1;ram[3][105]=0;ram[3][106]=1;ram[3][107]=1;ram[3][108]=0;ram[3][109]=1;ram[3][110]=1;ram[3][111]=0;ram[3][112]=0;ram[3][113]=1;ram[3][114]=1;ram[3][115]=0;ram[3][116]=1;ram[3][117]=1;ram[3][118]=1;ram[3][119]=1;ram[3][120]=1;ram[3][121]=1;ram[3][122]=0;ram[3][123]=1;ram[3][124]=1;ram[3][125]=0;ram[3][126]=0;ram[3][127]=1;ram[3][128]=0;ram[3][129]=1;ram[3][130]=1;ram[3][131]=0;ram[3][132]=1;ram[3][133]=1;ram[3][134]=1;ram[3][135]=0;ram[3][136]=0;
        ram[4][0]=1;ram[4][1]=1;ram[4][2]=1;ram[4][3]=1;ram[4][4]=1;ram[4][5]=1;ram[4][6]=0;ram[4][7]=0;ram[4][8]=0;ram[4][9]=0;ram[4][10]=1;ram[4][11]=0;ram[4][12]=1;ram[4][13]=1;ram[4][14]=1;ram[4][15]=0;ram[4][16]=1;ram[4][17]=0;ram[4][18]=1;ram[4][19]=1;ram[4][20]=1;ram[4][21]=1;ram[4][22]=0;ram[4][23]=1;ram[4][24]=0;ram[4][25]=1;ram[4][26]=1;ram[4][27]=1;ram[4][28]=1;ram[4][29]=0;ram[4][30]=0;ram[4][31]=1;ram[4][32]=1;ram[4][33]=1;ram[4][34]=1;ram[4][35]=0;ram[4][36]=1;ram[4][37]=1;ram[4][38]=0;ram[4][39]=0;ram[4][40]=0;ram[4][41]=1;ram[4][42]=0;ram[4][43]=1;ram[4][44]=1;ram[4][45]=1;ram[4][46]=0;ram[4][47]=1;ram[4][48]=1;ram[4][49]=0;ram[4][50]=0;ram[4][51]=1;ram[4][52]=1;ram[4][53]=1;ram[4][54]=1;ram[4][55]=1;ram[4][56]=1;ram[4][57]=1;ram[4][58]=1;ram[4][59]=0;ram[4][60]=1;ram[4][61]=1;ram[4][62]=0;ram[4][63]=1;ram[4][64]=1;ram[4][65]=1;ram[4][66]=1;ram[4][67]=1;ram[4][68]=0;ram[4][69]=0;ram[4][70]=0;ram[4][71]=1;ram[4][72]=0;ram[4][73]=0;ram[4][74]=0;ram[4][75]=1;ram[4][76]=1;ram[4][77]=1;ram[4][78]=1;ram[4][79]=1;ram[4][80]=1;ram[4][81]=1;ram[4][82]=0;ram[4][83]=1;ram[4][84]=1;ram[4][85]=0;ram[4][86]=0;ram[4][87]=1;ram[4][88]=1;ram[4][89]=1;ram[4][90]=0;ram[4][91]=1;ram[4][92]=1;ram[4][93]=0;ram[4][94]=1;ram[4][95]=1;ram[4][96]=0;ram[4][97]=0;ram[4][98]=0;ram[4][99]=1;ram[4][100]=0;ram[4][101]=0;ram[4][102]=1;ram[4][103]=1;ram[4][104]=0;ram[4][105]=1;ram[4][106]=1;ram[4][107]=1;ram[4][108]=1;ram[4][109]=1;ram[4][110]=0;ram[4][111]=0;ram[4][112]=1;ram[4][113]=1;ram[4][114]=0;ram[4][115]=1;ram[4][116]=0;ram[4][117]=0;ram[4][118]=0;ram[4][119]=1;ram[4][120]=0;ram[4][121]=1;ram[4][122]=1;ram[4][123]=1;ram[4][124]=1;ram[4][125]=0;ram[4][126]=0;ram[4][127]=1;ram[4][128]=0;ram[4][129]=1;ram[4][130]=1;ram[4][131]=0;ram[4][132]=0;ram[4][133]=1;ram[4][134]=1;ram[4][135]=0;ram[4][136]=1;
        ram[5][0]=1;ram[5][1]=0;ram[5][2]=1;ram[5][3]=0;ram[5][4]=0;ram[5][5]=1;ram[5][6]=0;ram[5][7]=1;ram[5][8]=0;ram[5][9]=1;ram[5][10]=1;ram[5][11]=0;ram[5][12]=1;ram[5][13]=0;ram[5][14]=0;ram[5][15]=1;ram[5][16]=1;ram[5][17]=0;ram[5][18]=0;ram[5][19]=1;ram[5][20]=1;ram[5][21]=1;ram[5][22]=1;ram[5][23]=1;ram[5][24]=1;ram[5][25]=0;ram[5][26]=1;ram[5][27]=1;ram[5][28]=0;ram[5][29]=1;ram[5][30]=1;ram[5][31]=1;ram[5][32]=1;ram[5][33]=1;ram[5][34]=1;ram[5][35]=0;ram[5][36]=1;ram[5][37]=1;ram[5][38]=0;ram[5][39]=0;ram[5][40]=1;ram[5][41]=1;ram[5][42]=1;ram[5][43]=1;ram[5][44]=0;ram[5][45]=0;ram[5][46]=1;ram[5][47]=1;ram[5][48]=0;ram[5][49]=1;ram[5][50]=0;ram[5][51]=1;ram[5][52]=1;ram[5][53]=0;ram[5][54]=0;ram[5][55]=0;ram[5][56]=1;ram[5][57]=1;ram[5][58]=1;ram[5][59]=1;ram[5][60]=1;ram[5][61]=1;ram[5][62]=1;ram[5][63]=1;ram[5][64]=0;ram[5][65]=1;ram[5][66]=1;ram[5][67]=1;ram[5][68]=0;ram[5][69]=0;ram[5][70]=1;ram[5][71]=1;ram[5][72]=1;ram[5][73]=1;ram[5][74]=1;ram[5][75]=1;ram[5][76]=0;ram[5][77]=1;ram[5][78]=1;ram[5][79]=0;ram[5][80]=1;ram[5][81]=0;ram[5][82]=0;ram[5][83]=1;ram[5][84]=1;ram[5][85]=0;ram[5][86]=0;ram[5][87]=0;ram[5][88]=1;ram[5][89]=1;ram[5][90]=0;ram[5][91]=1;ram[5][92]=0;ram[5][93]=1;ram[5][94]=0;ram[5][95]=0;ram[5][96]=0;ram[5][97]=1;ram[5][98]=0;ram[5][99]=1;ram[5][100]=0;ram[5][101]=0;ram[5][102]=0;ram[5][103]=1;ram[5][104]=1;ram[5][105]=1;ram[5][106]=1;ram[5][107]=1;ram[5][108]=1;ram[5][109]=1;ram[5][110]=1;ram[5][111]=1;ram[5][112]=0;ram[5][113]=1;ram[5][114]=0;ram[5][115]=0;ram[5][116]=0;ram[5][117]=1;ram[5][118]=0;ram[5][119]=0;ram[5][120]=0;ram[5][121]=1;ram[5][122]=1;ram[5][123]=1;ram[5][124]=1;ram[5][125]=0;ram[5][126]=1;ram[5][127]=1;ram[5][128]=1;ram[5][129]=1;ram[5][130]=0;ram[5][131]=1;ram[5][132]=1;ram[5][133]=1;ram[5][134]=1;ram[5][135]=0;ram[5][136]=0;
        ram[6][0]=1;ram[6][1]=1;ram[6][2]=0;ram[6][3]=0;ram[6][4]=0;ram[6][5]=1;ram[6][6]=1;ram[6][7]=1;ram[6][8]=1;ram[6][9]=1;ram[6][10]=1;ram[6][11]=0;ram[6][12]=1;ram[6][13]=0;ram[6][14]=0;ram[6][15]=1;ram[6][16]=0;ram[6][17]=1;ram[6][18]=1;ram[6][19]=0;ram[6][20]=0;ram[6][21]=1;ram[6][22]=1;ram[6][23]=0;ram[6][24]=0;ram[6][25]=1;ram[6][26]=0;ram[6][27]=1;ram[6][28]=0;ram[6][29]=1;ram[6][30]=1;ram[6][31]=1;ram[6][32]=0;ram[6][33]=0;ram[6][34]=1;ram[6][35]=0;ram[6][36]=1;ram[6][37]=0;ram[6][38]=1;ram[6][39]=1;ram[6][40]=1;ram[6][41]=1;ram[6][42]=0;ram[6][43]=1;ram[6][44]=1;ram[6][45]=1;ram[6][46]=0;ram[6][47]=1;ram[6][48]=1;ram[6][49]=1;ram[6][50]=1;ram[6][51]=1;ram[6][52]=1;ram[6][53]=1;ram[6][54]=0;ram[6][55]=0;ram[6][56]=0;ram[6][57]=1;ram[6][58]=0;ram[6][59]=1;ram[6][60]=0;ram[6][61]=1;ram[6][62]=1;ram[6][63]=1;ram[6][64]=1;ram[6][65]=1;ram[6][66]=1;ram[6][67]=0;ram[6][68]=1;ram[6][69]=1;ram[6][70]=1;ram[6][71]=0;ram[6][72]=0;ram[6][73]=0;ram[6][74]=1;ram[6][75]=1;ram[6][76]=1;ram[6][77]=1;ram[6][78]=1;ram[6][79]=0;ram[6][80]=1;ram[6][81]=1;ram[6][82]=0;ram[6][83]=0;ram[6][84]=1;ram[6][85]=0;ram[6][86]=0;ram[6][87]=1;ram[6][88]=1;ram[6][89]=1;ram[6][90]=1;ram[6][91]=0;ram[6][92]=1;ram[6][93]=1;ram[6][94]=0;ram[6][95]=0;ram[6][96]=1;ram[6][97]=1;ram[6][98]=1;ram[6][99]=1;ram[6][100]=1;ram[6][101]=1;ram[6][102]=1;ram[6][103]=1;ram[6][104]=0;ram[6][105]=0;ram[6][106]=0;ram[6][107]=1;ram[6][108]=0;ram[6][109]=1;ram[6][110]=0;ram[6][111]=1;ram[6][112]=0;ram[6][113]=0;ram[6][114]=0;ram[6][115]=1;ram[6][116]=1;ram[6][117]=1;ram[6][118]=1;ram[6][119]=0;ram[6][120]=0;ram[6][121]=1;ram[6][122]=1;ram[6][123]=0;ram[6][124]=1;ram[6][125]=1;ram[6][126]=1;ram[6][127]=1;ram[6][128]=0;ram[6][129]=1;ram[6][130]=1;ram[6][131]=1;ram[6][132]=1;ram[6][133]=1;ram[6][134]=1;ram[6][135]=1;ram[6][136]=1;
        ram[7][0]=1;ram[7][1]=1;ram[7][2]=1;ram[7][3]=1;ram[7][4]=0;ram[7][5]=1;ram[7][6]=1;ram[7][7]=1;ram[7][8]=1;ram[7][9]=0;ram[7][10]=1;ram[7][11]=1;ram[7][12]=0;ram[7][13]=1;ram[7][14]=0;ram[7][15]=1;ram[7][16]=1;ram[7][17]=1;ram[7][18]=1;ram[7][19]=1;ram[7][20]=1;ram[7][21]=1;ram[7][22]=1;ram[7][23]=0;ram[7][24]=0;ram[7][25]=1;ram[7][26]=0;ram[7][27]=0;ram[7][28]=1;ram[7][29]=1;ram[7][30]=1;ram[7][31]=1;ram[7][32]=0;ram[7][33]=0;ram[7][34]=0;ram[7][35]=1;ram[7][36]=1;ram[7][37]=1;ram[7][38]=1;ram[7][39]=1;ram[7][40]=0;ram[7][41]=0;ram[7][42]=1;ram[7][43]=1;ram[7][44]=1;ram[7][45]=1;ram[7][46]=0;ram[7][47]=1;ram[7][48]=0;ram[7][49]=0;ram[7][50]=1;ram[7][51]=0;ram[7][52]=0;ram[7][53]=0;ram[7][54]=0;ram[7][55]=1;ram[7][56]=1;ram[7][57]=1;ram[7][58]=1;ram[7][59]=1;ram[7][60]=1;ram[7][61]=1;ram[7][62]=1;ram[7][63]=0;ram[7][64]=1;ram[7][65]=0;ram[7][66]=1;ram[7][67]=0;ram[7][68]=0;ram[7][69]=1;ram[7][70]=1;ram[7][71]=0;ram[7][72]=0;ram[7][73]=0;ram[7][74]=1;ram[7][75]=1;ram[7][76]=0;ram[7][77]=0;ram[7][78]=1;ram[7][79]=1;ram[7][80]=1;ram[7][81]=1;ram[7][82]=1;ram[7][83]=0;ram[7][84]=1;ram[7][85]=0;ram[7][86]=1;ram[7][87]=0;ram[7][88]=0;ram[7][89]=0;ram[7][90]=1;ram[7][91]=1;ram[7][92]=1;ram[7][93]=0;ram[7][94]=1;ram[7][95]=1;ram[7][96]=1;ram[7][97]=1;ram[7][98]=1;ram[7][99]=1;ram[7][100]=1;ram[7][101]=1;ram[7][102]=1;ram[7][103]=1;ram[7][104]=1;ram[7][105]=0;ram[7][106]=1;ram[7][107]=0;ram[7][108]=1;ram[7][109]=0;ram[7][110]=0;ram[7][111]=1;ram[7][112]=0;ram[7][113]=1;ram[7][114]=1;ram[7][115]=1;ram[7][116]=0;ram[7][117]=0;ram[7][118]=1;ram[7][119]=1;ram[7][120]=0;ram[7][121]=1;ram[7][122]=1;ram[7][123]=0;ram[7][124]=0;ram[7][125]=1;ram[7][126]=1;ram[7][127]=1;ram[7][128]=1;ram[7][129]=1;ram[7][130]=1;ram[7][131]=1;ram[7][132]=1;ram[7][133]=0;ram[7][134]=0;ram[7][135]=1;ram[7][136]=0;
        ram[8][0]=1;ram[8][1]=1;ram[8][2]=0;ram[8][3]=1;ram[8][4]=0;ram[8][5]=0;ram[8][6]=1;ram[8][7]=1;ram[8][8]=0;ram[8][9]=1;ram[8][10]=1;ram[8][11]=1;ram[8][12]=1;ram[8][13]=1;ram[8][14]=1;ram[8][15]=0;ram[8][16]=0;ram[8][17]=1;ram[8][18]=0;ram[8][19]=1;ram[8][20]=1;ram[8][21]=1;ram[8][22]=1;ram[8][23]=1;ram[8][24]=1;ram[8][25]=0;ram[8][26]=0;ram[8][27]=1;ram[8][28]=1;ram[8][29]=0;ram[8][30]=1;ram[8][31]=1;ram[8][32]=0;ram[8][33]=1;ram[8][34]=1;ram[8][35]=1;ram[8][36]=0;ram[8][37]=1;ram[8][38]=0;ram[8][39]=1;ram[8][40]=0;ram[8][41]=1;ram[8][42]=1;ram[8][43]=0;ram[8][44]=0;ram[8][45]=1;ram[8][46]=1;ram[8][47]=1;ram[8][48]=0;ram[8][49]=1;ram[8][50]=0;ram[8][51]=1;ram[8][52]=1;ram[8][53]=1;ram[8][54]=1;ram[8][55]=1;ram[8][56]=1;ram[8][57]=0;ram[8][58]=1;ram[8][59]=1;ram[8][60]=1;ram[8][61]=1;ram[8][62]=0;ram[8][63]=0;ram[8][64]=1;ram[8][65]=1;ram[8][66]=1;ram[8][67]=1;ram[8][68]=1;ram[8][69]=1;ram[8][70]=1;ram[8][71]=1;ram[8][72]=1;ram[8][73]=1;ram[8][74]=1;ram[8][75]=1;ram[8][76]=1;ram[8][77]=1;ram[8][78]=1;ram[8][79]=0;ram[8][80]=0;ram[8][81]=1;ram[8][82]=1;ram[8][83]=1;ram[8][84]=0;ram[8][85]=1;ram[8][86]=0;ram[8][87]=1;ram[8][88]=1;ram[8][89]=1;ram[8][90]=1;ram[8][91]=0;ram[8][92]=0;ram[8][93]=1;ram[8][94]=0;ram[8][95]=0;ram[8][96]=0;ram[8][97]=1;ram[8][98]=1;ram[8][99]=1;ram[8][100]=1;ram[8][101]=1;ram[8][102]=1;ram[8][103]=1;ram[8][104]=1;ram[8][105]=1;ram[8][106]=1;ram[8][107]=1;ram[8][108]=1;ram[8][109]=0;ram[8][110]=1;ram[8][111]=0;ram[8][112]=0;ram[8][113]=0;ram[8][114]=1;ram[8][115]=1;ram[8][116]=0;ram[8][117]=0;ram[8][118]=1;ram[8][119]=1;ram[8][120]=0;ram[8][121]=1;ram[8][122]=1;ram[8][123]=1;ram[8][124]=0;ram[8][125]=0;ram[8][126]=1;ram[8][127]=0;ram[8][128]=1;ram[8][129]=1;ram[8][130]=1;ram[8][131]=1;ram[8][132]=0;ram[8][133]=1;ram[8][134]=1;ram[8][135]=0;ram[8][136]=1;
        ram[9][0]=1;ram[9][1]=0;ram[9][2]=1;ram[9][3]=1;ram[9][4]=1;ram[9][5]=0;ram[9][6]=1;ram[9][7]=1;ram[9][8]=0;ram[9][9]=1;ram[9][10]=0;ram[9][11]=1;ram[9][12]=1;ram[9][13]=0;ram[9][14]=1;ram[9][15]=0;ram[9][16]=1;ram[9][17]=1;ram[9][18]=1;ram[9][19]=1;ram[9][20]=1;ram[9][21]=1;ram[9][22]=0;ram[9][23]=1;ram[9][24]=1;ram[9][25]=1;ram[9][26]=1;ram[9][27]=0;ram[9][28]=1;ram[9][29]=0;ram[9][30]=0;ram[9][31]=0;ram[9][32]=0;ram[9][33]=1;ram[9][34]=1;ram[9][35]=1;ram[9][36]=0;ram[9][37]=1;ram[9][38]=1;ram[9][39]=0;ram[9][40]=1;ram[9][41]=1;ram[9][42]=1;ram[9][43]=1;ram[9][44]=1;ram[9][45]=0;ram[9][46]=1;ram[9][47]=1;ram[9][48]=1;ram[9][49]=0;ram[9][50]=1;ram[9][51]=0;ram[9][52]=1;ram[9][53]=1;ram[9][54]=0;ram[9][55]=0;ram[9][56]=0;ram[9][57]=1;ram[9][58]=1;ram[9][59]=0;ram[9][60]=1;ram[9][61]=1;ram[9][62]=1;ram[9][63]=0;ram[9][64]=1;ram[9][65]=1;ram[9][66]=1;ram[9][67]=1;ram[9][68]=1;ram[9][69]=0;ram[9][70]=1;ram[9][71]=1;ram[9][72]=1;ram[9][73]=1;ram[9][74]=0;ram[9][75]=1;ram[9][76]=0;ram[9][77]=1;ram[9][78]=0;ram[9][79]=1;ram[9][80]=1;ram[9][81]=1;ram[9][82]=1;ram[9][83]=1;ram[9][84]=0;ram[9][85]=0;ram[9][86]=0;ram[9][87]=1;ram[9][88]=1;ram[9][89]=0;ram[9][90]=0;ram[9][91]=0;ram[9][92]=1;ram[9][93]=1;ram[9][94]=0;ram[9][95]=1;ram[9][96]=0;ram[9][97]=1;ram[9][98]=0;ram[9][99]=1;ram[9][100]=0;ram[9][101]=1;ram[9][102]=1;ram[9][103]=1;ram[9][104]=1;ram[9][105]=1;ram[9][106]=0;ram[9][107]=1;ram[9][108]=1;ram[9][109]=1;ram[9][110]=1;ram[9][111]=0;ram[9][112]=1;ram[9][113]=1;ram[9][114]=1;ram[9][115]=0;ram[9][116]=1;ram[9][117]=1;ram[9][118]=1;ram[9][119]=0;ram[9][120]=0;ram[9][121]=1;ram[9][122]=0;ram[9][123]=0;ram[9][124]=0;ram[9][125]=1;ram[9][126]=1;ram[9][127]=1;ram[9][128]=1;ram[9][129]=1;ram[9][130]=1;ram[9][131]=0;ram[9][132]=1;ram[9][133]=0;ram[9][134]=1;ram[9][135]=1;ram[9][136]=1;
        ram[10][0]=1;ram[10][1]=1;ram[10][2]=1;ram[10][3]=1;ram[10][4]=0;ram[10][5]=1;ram[10][6]=1;ram[10][7]=1;ram[10][8]=1;ram[10][9]=1;ram[10][10]=1;ram[10][11]=1;ram[10][12]=1;ram[10][13]=1;ram[10][14]=1;ram[10][15]=1;ram[10][16]=1;ram[10][17]=0;ram[10][18]=1;ram[10][19]=1;ram[10][20]=1;ram[10][21]=1;ram[10][22]=1;ram[10][23]=1;ram[10][24]=1;ram[10][25]=1;ram[10][26]=0;ram[10][27]=0;ram[10][28]=0;ram[10][29]=1;ram[10][30]=1;ram[10][31]=1;ram[10][32]=0;ram[10][33]=0;ram[10][34]=1;ram[10][35]=1;ram[10][36]=0;ram[10][37]=1;ram[10][38]=0;ram[10][39]=1;ram[10][40]=0;ram[10][41]=1;ram[10][42]=1;ram[10][43]=0;ram[10][44]=1;ram[10][45]=0;ram[10][46]=0;ram[10][47]=1;ram[10][48]=0;ram[10][49]=1;ram[10][50]=1;ram[10][51]=1;ram[10][52]=1;ram[10][53]=1;ram[10][54]=0;ram[10][55]=1;ram[10][56]=1;ram[10][57]=0;ram[10][58]=0;ram[10][59]=0;ram[10][60]=1;ram[10][61]=1;ram[10][62]=1;ram[10][63]=0;ram[10][64]=0;ram[10][65]=0;ram[10][66]=0;ram[10][67]=1;ram[10][68]=0;ram[10][69]=0;ram[10][70]=1;ram[10][71]=1;ram[10][72]=1;ram[10][73]=1;ram[10][74]=1;ram[10][75]=1;ram[10][76]=1;ram[10][77]=1;ram[10][78]=1;ram[10][79]=0;ram[10][80]=1;ram[10][81]=0;ram[10][82]=1;ram[10][83]=1;ram[10][84]=1;ram[10][85]=0;ram[10][86]=1;ram[10][87]=0;ram[10][88]=1;ram[10][89]=0;ram[10][90]=0;ram[10][91]=1;ram[10][92]=0;ram[10][93]=1;ram[10][94]=0;ram[10][95]=1;ram[10][96]=1;ram[10][97]=0;ram[10][98]=1;ram[10][99]=1;ram[10][100]=1;ram[10][101]=1;ram[10][102]=0;ram[10][103]=0;ram[10][104]=1;ram[10][105]=1;ram[10][106]=0;ram[10][107]=0;ram[10][108]=0;ram[10][109]=0;ram[10][110]=1;ram[10][111]=1;ram[10][112]=1;ram[10][113]=1;ram[10][114]=1;ram[10][115]=1;ram[10][116]=1;ram[10][117]=0;ram[10][118]=1;ram[10][119]=1;ram[10][120]=1;ram[10][121]=1;ram[10][122]=1;ram[10][123]=1;ram[10][124]=0;ram[10][125]=1;ram[10][126]=0;ram[10][127]=1;ram[10][128]=1;ram[10][129]=1;ram[10][130]=1;ram[10][131]=1;ram[10][132]=1;ram[10][133]=1;ram[10][134]=1;ram[10][135]=1;ram[10][136]=0;
        ram[11][0]=1;ram[11][1]=1;ram[11][2]=1;ram[11][3]=1;ram[11][4]=1;ram[11][5]=1;ram[11][6]=1;ram[11][7]=0;ram[11][8]=1;ram[11][9]=0;ram[11][10]=1;ram[11][11]=1;ram[11][12]=1;ram[11][13]=1;ram[11][14]=1;ram[11][15]=1;ram[11][16]=0;ram[11][17]=1;ram[11][18]=1;ram[11][19]=0;ram[11][20]=1;ram[11][21]=1;ram[11][22]=1;ram[11][23]=1;ram[11][24]=0;ram[11][25]=1;ram[11][26]=0;ram[11][27]=1;ram[11][28]=0;ram[11][29]=0;ram[11][30]=0;ram[11][31]=0;ram[11][32]=1;ram[11][33]=1;ram[11][34]=1;ram[11][35]=1;ram[11][36]=0;ram[11][37]=0;ram[11][38]=1;ram[11][39]=1;ram[11][40]=0;ram[11][41]=1;ram[11][42]=1;ram[11][43]=1;ram[11][44]=0;ram[11][45]=1;ram[11][46]=0;ram[11][47]=1;ram[11][48]=1;ram[11][49]=1;ram[11][50]=1;ram[11][51]=1;ram[11][52]=0;ram[11][53]=0;ram[11][54]=0;ram[11][55]=1;ram[11][56]=1;ram[11][57]=1;ram[11][58]=1;ram[11][59]=1;ram[11][60]=1;ram[11][61]=0;ram[11][62]=1;ram[11][63]=0;ram[11][64]=1;ram[11][65]=1;ram[11][66]=1;ram[11][67]=1;ram[11][68]=1;ram[11][69]=1;ram[11][70]=1;ram[11][71]=1;ram[11][72]=1;ram[11][73]=0;ram[11][74]=0;ram[11][75]=1;ram[11][76]=1;ram[11][77]=0;ram[11][78]=0;ram[11][79]=1;ram[11][80]=1;ram[11][81]=0;ram[11][82]=0;ram[11][83]=1;ram[11][84]=1;ram[11][85]=1;ram[11][86]=1;ram[11][87]=0;ram[11][88]=1;ram[11][89]=0;ram[11][90]=0;ram[11][91]=1;ram[11][92]=0;ram[11][93]=0;ram[11][94]=0;ram[11][95]=1;ram[11][96]=1;ram[11][97]=1;ram[11][98]=1;ram[11][99]=0;ram[11][100]=0;ram[11][101]=0;ram[11][102]=0;ram[11][103]=0;ram[11][104]=1;ram[11][105]=0;ram[11][106]=1;ram[11][107]=1;ram[11][108]=1;ram[11][109]=0;ram[11][110]=1;ram[11][111]=0;ram[11][112]=1;ram[11][113]=1;ram[11][114]=1;ram[11][115]=0;ram[11][116]=1;ram[11][117]=1;ram[11][118]=1;ram[11][119]=1;ram[11][120]=1;ram[11][121]=0;ram[11][122]=1;ram[11][123]=1;ram[11][124]=0;ram[11][125]=0;ram[11][126]=1;ram[11][127]=0;ram[11][128]=1;ram[11][129]=0;ram[11][130]=0;ram[11][131]=0;ram[11][132]=1;ram[11][133]=0;ram[11][134]=0;ram[11][135]=0;ram[11][136]=1;
        ram[12][0]=0;ram[12][1]=0;ram[12][2]=1;ram[12][3]=1;ram[12][4]=0;ram[12][5]=0;ram[12][6]=1;ram[12][7]=0;ram[12][8]=1;ram[12][9]=0;ram[12][10]=0;ram[12][11]=0;ram[12][12]=0;ram[12][13]=1;ram[12][14]=1;ram[12][15]=0;ram[12][16]=1;ram[12][17]=1;ram[12][18]=1;ram[12][19]=0;ram[12][20]=0;ram[12][21]=1;ram[12][22]=1;ram[12][23]=1;ram[12][24]=1;ram[12][25]=1;ram[12][26]=0;ram[12][27]=1;ram[12][28]=1;ram[12][29]=1;ram[12][30]=1;ram[12][31]=0;ram[12][32]=0;ram[12][33]=1;ram[12][34]=1;ram[12][35]=1;ram[12][36]=1;ram[12][37]=0;ram[12][38]=1;ram[12][39]=0;ram[12][40]=1;ram[12][41]=0;ram[12][42]=1;ram[12][43]=1;ram[12][44]=1;ram[12][45]=0;ram[12][46]=0;ram[12][47]=0;ram[12][48]=1;ram[12][49]=1;ram[12][50]=1;ram[12][51]=0;ram[12][52]=1;ram[12][53]=1;ram[12][54]=0;ram[12][55]=1;ram[12][56]=0;ram[12][57]=1;ram[12][58]=1;ram[12][59]=1;ram[12][60]=0;ram[12][61]=0;ram[12][62]=0;ram[12][63]=1;ram[12][64]=1;ram[12][65]=1;ram[12][66]=1;ram[12][67]=1;ram[12][68]=0;ram[12][69]=0;ram[12][70]=1;ram[12][71]=0;ram[12][72]=1;ram[12][73]=0;ram[12][74]=0;ram[12][75]=0;ram[12][76]=0;ram[12][77]=0;ram[12][78]=0;ram[12][79]=0;ram[12][80]=1;ram[12][81]=1;ram[12][82]=0;ram[12][83]=0;ram[12][84]=1;ram[12][85]=1;ram[12][86]=0;ram[12][87]=1;ram[12][88]=0;ram[12][89]=1;ram[12][90]=1;ram[12][91]=1;ram[12][92]=1;ram[12][93]=1;ram[12][94]=1;ram[12][95]=0;ram[12][96]=1;ram[12][97]=1;ram[12][98]=1;ram[12][99]=1;ram[12][100]=1;ram[12][101]=1;ram[12][102]=1;ram[12][103]=0;ram[12][104]=1;ram[12][105]=1;ram[12][106]=0;ram[12][107]=1;ram[12][108]=1;ram[12][109]=0;ram[12][110]=1;ram[12][111]=0;ram[12][112]=0;ram[12][113]=1;ram[12][114]=1;ram[12][115]=1;ram[12][116]=0;ram[12][117]=1;ram[12][118]=1;ram[12][119]=1;ram[12][120]=0;ram[12][121]=1;ram[12][122]=1;ram[12][123]=1;ram[12][124]=0;ram[12][125]=0;ram[12][126]=0;ram[12][127]=1;ram[12][128]=1;ram[12][129]=0;ram[12][130]=1;ram[12][131]=0;ram[12][132]=1;ram[12][133]=1;ram[12][134]=1;ram[12][135]=0;ram[12][136]=0;
        ram[13][0]=1;ram[13][1]=0;ram[13][2]=0;ram[13][3]=0;ram[13][4]=1;ram[13][5]=1;ram[13][6]=0;ram[13][7]=1;ram[13][8]=1;ram[13][9]=0;ram[13][10]=1;ram[13][11]=0;ram[13][12]=0;ram[13][13]=1;ram[13][14]=1;ram[13][15]=1;ram[13][16]=1;ram[13][17]=1;ram[13][18]=0;ram[13][19]=0;ram[13][20]=1;ram[13][21]=1;ram[13][22]=1;ram[13][23]=0;ram[13][24]=1;ram[13][25]=1;ram[13][26]=0;ram[13][27]=1;ram[13][28]=1;ram[13][29]=1;ram[13][30]=1;ram[13][31]=1;ram[13][32]=1;ram[13][33]=1;ram[13][34]=1;ram[13][35]=1;ram[13][36]=0;ram[13][37]=0;ram[13][38]=1;ram[13][39]=1;ram[13][40]=0;ram[13][41]=1;ram[13][42]=1;ram[13][43]=1;ram[13][44]=1;ram[13][45]=0;ram[13][46]=0;ram[13][47]=1;ram[13][48]=1;ram[13][49]=0;ram[13][50]=1;ram[13][51]=1;ram[13][52]=0;ram[13][53]=0;ram[13][54]=1;ram[13][55]=1;ram[13][56]=1;ram[13][57]=1;ram[13][58]=1;ram[13][59]=0;ram[13][60]=1;ram[13][61]=1;ram[13][62]=1;ram[13][63]=1;ram[13][64]=1;ram[13][65]=1;ram[13][66]=1;ram[13][67]=1;ram[13][68]=1;ram[13][69]=1;ram[13][70]=1;ram[13][71]=0;ram[13][72]=1;ram[13][73]=0;ram[13][74]=1;ram[13][75]=0;ram[13][76]=1;ram[13][77]=1;ram[13][78]=0;ram[13][79]=0;ram[13][80]=1;ram[13][81]=1;ram[13][82]=0;ram[13][83]=0;ram[13][84]=1;ram[13][85]=1;ram[13][86]=1;ram[13][87]=0;ram[13][88]=1;ram[13][89]=1;ram[13][90]=1;ram[13][91]=1;ram[13][92]=0;ram[13][93]=0;ram[13][94]=1;ram[13][95]=1;ram[13][96]=1;ram[13][97]=1;ram[13][98]=0;ram[13][99]=1;ram[13][100]=1;ram[13][101]=1;ram[13][102]=1;ram[13][103]=0;ram[13][104]=0;ram[13][105]=1;ram[13][106]=0;ram[13][107]=1;ram[13][108]=0;ram[13][109]=0;ram[13][110]=1;ram[13][111]=1;ram[13][112]=1;ram[13][113]=1;ram[13][114]=0;ram[13][115]=0;ram[13][116]=1;ram[13][117]=1;ram[13][118]=1;ram[13][119]=0;ram[13][120]=1;ram[13][121]=0;ram[13][122]=0;ram[13][123]=1;ram[13][124]=1;ram[13][125]=0;ram[13][126]=1;ram[13][127]=0;ram[13][128]=0;ram[13][129]=1;ram[13][130]=1;ram[13][131]=0;ram[13][132]=1;ram[13][133]=0;ram[13][134]=1;ram[13][135]=0;ram[13][136]=0;
        ram[14][0]=1;ram[14][1]=0;ram[14][2]=1;ram[14][3]=1;ram[14][4]=1;ram[14][5]=1;ram[14][6]=0;ram[14][7]=1;ram[14][8]=0;ram[14][9]=0;ram[14][10]=1;ram[14][11]=1;ram[14][12]=1;ram[14][13]=1;ram[14][14]=1;ram[14][15]=1;ram[14][16]=0;ram[14][17]=1;ram[14][18]=0;ram[14][19]=1;ram[14][20]=1;ram[14][21]=1;ram[14][22]=1;ram[14][23]=1;ram[14][24]=1;ram[14][25]=1;ram[14][26]=1;ram[14][27]=0;ram[14][28]=0;ram[14][29]=0;ram[14][30]=1;ram[14][31]=1;ram[14][32]=1;ram[14][33]=1;ram[14][34]=1;ram[14][35]=1;ram[14][36]=0;ram[14][37]=1;ram[14][38]=1;ram[14][39]=1;ram[14][40]=1;ram[14][41]=1;ram[14][42]=1;ram[14][43]=1;ram[14][44]=1;ram[14][45]=1;ram[14][46]=1;ram[14][47]=1;ram[14][48]=1;ram[14][49]=1;ram[14][50]=1;ram[14][51]=1;ram[14][52]=0;ram[14][53]=1;ram[14][54]=0;ram[14][55]=0;ram[14][56]=0;ram[14][57]=1;ram[14][58]=1;ram[14][59]=1;ram[14][60]=0;ram[14][61]=1;ram[14][62]=0;ram[14][63]=1;ram[14][64]=1;ram[14][65]=1;ram[14][66]=1;ram[14][67]=1;ram[14][68]=1;ram[14][69]=1;ram[14][70]=1;ram[14][71]=1;ram[14][72]=0;ram[14][73]=1;ram[14][74]=1;ram[14][75]=0;ram[14][76]=1;ram[14][77]=1;ram[14][78]=1;ram[14][79]=0;ram[14][80]=0;ram[14][81]=1;ram[14][82]=1;ram[14][83]=1;ram[14][84]=1;ram[14][85]=1;ram[14][86]=1;ram[14][87]=1;ram[14][88]=1;ram[14][89]=0;ram[14][90]=0;ram[14][91]=0;ram[14][92]=0;ram[14][93]=0;ram[14][94]=0;ram[14][95]=1;ram[14][96]=1;ram[14][97]=1;ram[14][98]=1;ram[14][99]=0;ram[14][100]=0;ram[14][101]=1;ram[14][102]=1;ram[14][103]=1;ram[14][104]=1;ram[14][105]=0;ram[14][106]=1;ram[14][107]=1;ram[14][108]=1;ram[14][109]=1;ram[14][110]=1;ram[14][111]=1;ram[14][112]=1;ram[14][113]=0;ram[14][114]=1;ram[14][115]=1;ram[14][116]=1;ram[14][117]=1;ram[14][118]=1;ram[14][119]=1;ram[14][120]=1;ram[14][121]=1;ram[14][122]=1;ram[14][123]=1;ram[14][124]=1;ram[14][125]=0;ram[14][126]=0;ram[14][127]=1;ram[14][128]=0;ram[14][129]=1;ram[14][130]=1;ram[14][131]=0;ram[14][132]=0;ram[14][133]=0;ram[14][134]=1;ram[14][135]=0;ram[14][136]=1;
        ram[15][0]=1;ram[15][1]=1;ram[15][2]=0;ram[15][3]=1;ram[15][4]=1;ram[15][5]=1;ram[15][6]=1;ram[15][7]=0;ram[15][8]=1;ram[15][9]=0;ram[15][10]=1;ram[15][11]=1;ram[15][12]=1;ram[15][13]=1;ram[15][14]=1;ram[15][15]=1;ram[15][16]=0;ram[15][17]=1;ram[15][18]=0;ram[15][19]=1;ram[15][20]=0;ram[15][21]=1;ram[15][22]=0;ram[15][23]=0;ram[15][24]=1;ram[15][25]=0;ram[15][26]=0;ram[15][27]=1;ram[15][28]=1;ram[15][29]=1;ram[15][30]=1;ram[15][31]=1;ram[15][32]=1;ram[15][33]=1;ram[15][34]=1;ram[15][35]=1;ram[15][36]=0;ram[15][37]=1;ram[15][38]=1;ram[15][39]=1;ram[15][40]=1;ram[15][41]=1;ram[15][42]=1;ram[15][43]=0;ram[15][44]=1;ram[15][45]=0;ram[15][46]=1;ram[15][47]=1;ram[15][48]=0;ram[15][49]=0;ram[15][50]=1;ram[15][51]=1;ram[15][52]=0;ram[15][53]=1;ram[15][54]=1;ram[15][55]=1;ram[15][56]=1;ram[15][57]=1;ram[15][58]=0;ram[15][59]=0;ram[15][60]=1;ram[15][61]=1;ram[15][62]=1;ram[15][63]=1;ram[15][64]=1;ram[15][65]=1;ram[15][66]=1;ram[15][67]=0;ram[15][68]=0;ram[15][69]=1;ram[15][70]=1;ram[15][71]=0;ram[15][72]=1;ram[15][73]=1;ram[15][74]=1;ram[15][75]=1;ram[15][76]=1;ram[15][77]=1;ram[15][78]=0;ram[15][79]=0;ram[15][80]=0;ram[15][81]=1;ram[15][82]=1;ram[15][83]=1;ram[15][84]=0;ram[15][85]=1;ram[15][86]=1;ram[15][87]=0;ram[15][88]=1;ram[15][89]=1;ram[15][90]=1;ram[15][91]=1;ram[15][92]=0;ram[15][93]=0;ram[15][94]=1;ram[15][95]=0;ram[15][96]=1;ram[15][97]=1;ram[15][98]=0;ram[15][99]=1;ram[15][100]=0;ram[15][101]=1;ram[15][102]=1;ram[15][103]=1;ram[15][104]=0;ram[15][105]=1;ram[15][106]=1;ram[15][107]=1;ram[15][108]=1;ram[15][109]=1;ram[15][110]=1;ram[15][111]=1;ram[15][112]=0;ram[15][113]=0;ram[15][114]=1;ram[15][115]=1;ram[15][116]=1;ram[15][117]=1;ram[15][118]=0;ram[15][119]=1;ram[15][120]=0;ram[15][121]=1;ram[15][122]=1;ram[15][123]=1;ram[15][124]=1;ram[15][125]=1;ram[15][126]=1;ram[15][127]=1;ram[15][128]=1;ram[15][129]=0;ram[15][130]=0;ram[15][131]=0;ram[15][132]=1;ram[15][133]=1;ram[15][134]=1;ram[15][135]=0;ram[15][136]=0;
        ram[16][0]=1;ram[16][1]=0;ram[16][2]=1;ram[16][3]=0;ram[16][4]=1;ram[16][5]=0;ram[16][6]=0;ram[16][7]=1;ram[16][8]=1;ram[16][9]=0;ram[16][10]=0;ram[16][11]=0;ram[16][12]=1;ram[16][13]=1;ram[16][14]=1;ram[16][15]=1;ram[16][16]=0;ram[16][17]=1;ram[16][18]=0;ram[16][19]=0;ram[16][20]=1;ram[16][21]=1;ram[16][22]=1;ram[16][23]=1;ram[16][24]=0;ram[16][25]=1;ram[16][26]=1;ram[16][27]=1;ram[16][28]=0;ram[16][29]=0;ram[16][30]=1;ram[16][31]=1;ram[16][32]=1;ram[16][33]=0;ram[16][34]=1;ram[16][35]=1;ram[16][36]=1;ram[16][37]=1;ram[16][38]=0;ram[16][39]=1;ram[16][40]=1;ram[16][41]=1;ram[16][42]=1;ram[16][43]=1;ram[16][44]=0;ram[16][45]=1;ram[16][46]=1;ram[16][47]=1;ram[16][48]=1;ram[16][49]=0;ram[16][50]=1;ram[16][51]=1;ram[16][52]=1;ram[16][53]=0;ram[16][54]=0;ram[16][55]=1;ram[16][56]=1;ram[16][57]=0;ram[16][58]=1;ram[16][59]=1;ram[16][60]=0;ram[16][61]=1;ram[16][62]=1;ram[16][63]=1;ram[16][64]=1;ram[16][65]=1;ram[16][66]=0;ram[16][67]=0;ram[16][68]=1;ram[16][69]=0;ram[16][70]=1;ram[16][71]=1;ram[16][72]=0;ram[16][73]=1;ram[16][74]=1;ram[16][75]=0;ram[16][76]=0;ram[16][77]=0;ram[16][78]=0;ram[16][79]=1;ram[16][80]=1;ram[16][81]=0;ram[16][82]=1;ram[16][83]=1;ram[16][84]=0;ram[16][85]=0;ram[16][86]=1;ram[16][87]=1;ram[16][88]=0;ram[16][89]=1;ram[16][90]=0;ram[16][91]=0;ram[16][92]=1;ram[16][93]=1;ram[16][94]=0;ram[16][95]=1;ram[16][96]=1;ram[16][97]=0;ram[16][98]=1;ram[16][99]=1;ram[16][100]=1;ram[16][101]=1;ram[16][102]=1;ram[16][103]=1;ram[16][104]=0;ram[16][105]=1;ram[16][106]=1;ram[16][107]=1;ram[16][108]=1;ram[16][109]=0;ram[16][110]=1;ram[16][111]=0;ram[16][112]=0;ram[16][113]=1;ram[16][114]=1;ram[16][115]=1;ram[16][116]=0;ram[16][117]=1;ram[16][118]=0;ram[16][119]=1;ram[16][120]=0;ram[16][121]=1;ram[16][122]=1;ram[16][123]=1;ram[16][124]=1;ram[16][125]=1;ram[16][126]=1;ram[16][127]=1;ram[16][128]=1;ram[16][129]=0;ram[16][130]=0;ram[16][131]=0;ram[16][132]=0;ram[16][133]=1;ram[16][134]=1;ram[16][135]=0;ram[16][136]=0;
        ram[17][0]=1;ram[17][1]=1;ram[17][2]=1;ram[17][3]=0;ram[17][4]=1;ram[17][5]=1;ram[17][6]=0;ram[17][7]=0;ram[17][8]=1;ram[17][9]=1;ram[17][10]=1;ram[17][11]=0;ram[17][12]=1;ram[17][13]=1;ram[17][14]=1;ram[17][15]=0;ram[17][16]=0;ram[17][17]=0;ram[17][18]=1;ram[17][19]=0;ram[17][20]=1;ram[17][21]=1;ram[17][22]=1;ram[17][23]=1;ram[17][24]=1;ram[17][25]=1;ram[17][26]=1;ram[17][27]=0;ram[17][28]=1;ram[17][29]=0;ram[17][30]=0;ram[17][31]=1;ram[17][32]=1;ram[17][33]=1;ram[17][34]=1;ram[17][35]=1;ram[17][36]=0;ram[17][37]=1;ram[17][38]=1;ram[17][39]=1;ram[17][40]=1;ram[17][41]=0;ram[17][42]=0;ram[17][43]=0;ram[17][44]=1;ram[17][45]=0;ram[17][46]=0;ram[17][47]=0;ram[17][48]=1;ram[17][49]=1;ram[17][50]=1;ram[17][51]=0;ram[17][52]=1;ram[17][53]=0;ram[17][54]=0;ram[17][55]=1;ram[17][56]=1;ram[17][57]=1;ram[17][58]=0;ram[17][59]=0;ram[17][60]=1;ram[17][61]=0;ram[17][62]=1;ram[17][63]=0;ram[17][64]=1;ram[17][65]=0;ram[17][66]=1;ram[17][67]=1;ram[17][68]=1;ram[17][69]=0;ram[17][70]=0;ram[17][71]=1;ram[17][72]=1;ram[17][73]=1;ram[17][74]=1;ram[17][75]=1;ram[17][76]=1;ram[17][77]=1;ram[17][78]=1;ram[17][79]=0;ram[17][80]=1;ram[17][81]=1;ram[17][82]=0;ram[17][83]=1;ram[17][84]=0;ram[17][85]=1;ram[17][86]=0;ram[17][87]=1;ram[17][88]=0;ram[17][89]=0;ram[17][90]=1;ram[17][91]=0;ram[17][92]=1;ram[17][93]=1;ram[17][94]=1;ram[17][95]=1;ram[17][96]=0;ram[17][97]=1;ram[17][98]=0;ram[17][99]=1;ram[17][100]=0;ram[17][101]=1;ram[17][102]=1;ram[17][103]=1;ram[17][104]=1;ram[17][105]=1;ram[17][106]=1;ram[17][107]=1;ram[17][108]=1;ram[17][109]=1;ram[17][110]=1;ram[17][111]=0;ram[17][112]=1;ram[17][113]=1;ram[17][114]=0;ram[17][115]=1;ram[17][116]=1;ram[17][117]=1;ram[17][118]=1;ram[17][119]=0;ram[17][120]=1;ram[17][121]=1;ram[17][122]=1;ram[17][123]=0;ram[17][124]=1;ram[17][125]=1;ram[17][126]=1;ram[17][127]=1;ram[17][128]=1;ram[17][129]=1;ram[17][130]=1;ram[17][131]=1;ram[17][132]=1;ram[17][133]=0;ram[17][134]=1;ram[17][135]=0;ram[17][136]=1;
        ram[18][0]=1;ram[18][1]=1;ram[18][2]=0;ram[18][3]=1;ram[18][4]=0;ram[18][5]=0;ram[18][6]=1;ram[18][7]=1;ram[18][8]=1;ram[18][9]=1;ram[18][10]=1;ram[18][11]=1;ram[18][12]=1;ram[18][13]=1;ram[18][14]=0;ram[18][15]=1;ram[18][16]=1;ram[18][17]=1;ram[18][18]=0;ram[18][19]=1;ram[18][20]=0;ram[18][21]=1;ram[18][22]=1;ram[18][23]=0;ram[18][24]=1;ram[18][25]=1;ram[18][26]=0;ram[18][27]=0;ram[18][28]=1;ram[18][29]=1;ram[18][30]=0;ram[18][31]=1;ram[18][32]=1;ram[18][33]=0;ram[18][34]=0;ram[18][35]=1;ram[18][36]=1;ram[18][37]=1;ram[18][38]=1;ram[18][39]=0;ram[18][40]=1;ram[18][41]=1;ram[18][42]=0;ram[18][43]=1;ram[18][44]=1;ram[18][45]=1;ram[18][46]=1;ram[18][47]=1;ram[18][48]=0;ram[18][49]=1;ram[18][50]=0;ram[18][51]=0;ram[18][52]=1;ram[18][53]=0;ram[18][54]=0;ram[18][55]=1;ram[18][56]=1;ram[18][57]=1;ram[18][58]=1;ram[18][59]=1;ram[18][60]=1;ram[18][61]=1;ram[18][62]=0;ram[18][63]=0;ram[18][64]=1;ram[18][65]=0;ram[18][66]=0;ram[18][67]=1;ram[18][68]=1;ram[18][69]=1;ram[18][70]=0;ram[18][71]=0;ram[18][72]=1;ram[18][73]=0;ram[18][74]=1;ram[18][75]=0;ram[18][76]=0;ram[18][77]=1;ram[18][78]=1;ram[18][79]=0;ram[18][80]=1;ram[18][81]=1;ram[18][82]=0;ram[18][83]=1;ram[18][84]=1;ram[18][85]=1;ram[18][86]=1;ram[18][87]=0;ram[18][88]=0;ram[18][89]=1;ram[18][90]=1;ram[18][91]=1;ram[18][92]=0;ram[18][93]=0;ram[18][94]=1;ram[18][95]=1;ram[18][96]=1;ram[18][97]=0;ram[18][98]=1;ram[18][99]=1;ram[18][100]=0;ram[18][101]=1;ram[18][102]=0;ram[18][103]=1;ram[18][104]=1;ram[18][105]=1;ram[18][106]=1;ram[18][107]=1;ram[18][108]=1;ram[18][109]=0;ram[18][110]=0;ram[18][111]=0;ram[18][112]=0;ram[18][113]=1;ram[18][114]=0;ram[18][115]=0;ram[18][116]=1;ram[18][117]=1;ram[18][118]=1;ram[18][119]=0;ram[18][120]=1;ram[18][121]=1;ram[18][122]=0;ram[18][123]=1;ram[18][124]=0;ram[18][125]=0;ram[18][126]=1;ram[18][127]=0;ram[18][128]=0;ram[18][129]=1;ram[18][130]=1;ram[18][131]=1;ram[18][132]=1;ram[18][133]=0;ram[18][134]=1;ram[18][135]=0;ram[18][136]=1;
        ram[19][0]=1;ram[19][1]=0;ram[19][2]=1;ram[19][3]=0;ram[19][4]=0;ram[19][5]=1;ram[19][6]=1;ram[19][7]=1;ram[19][8]=0;ram[19][9]=0;ram[19][10]=1;ram[19][11]=1;ram[19][12]=1;ram[19][13]=1;ram[19][14]=1;ram[19][15]=1;ram[19][16]=0;ram[19][17]=0;ram[19][18]=1;ram[19][19]=1;ram[19][20]=1;ram[19][21]=0;ram[19][22]=1;ram[19][23]=1;ram[19][24]=1;ram[19][25]=1;ram[19][26]=0;ram[19][27]=1;ram[19][28]=0;ram[19][29]=0;ram[19][30]=1;ram[19][31]=1;ram[19][32]=1;ram[19][33]=0;ram[19][34]=1;ram[19][35]=0;ram[19][36]=1;ram[19][37]=0;ram[19][38]=1;ram[19][39]=1;ram[19][40]=0;ram[19][41]=1;ram[19][42]=0;ram[19][43]=1;ram[19][44]=0;ram[19][45]=1;ram[19][46]=1;ram[19][47]=1;ram[19][48]=1;ram[19][49]=0;ram[19][50]=1;ram[19][51]=1;ram[19][52]=0;ram[19][53]=0;ram[19][54]=0;ram[19][55]=0;ram[19][56]=1;ram[19][57]=0;ram[19][58]=1;ram[19][59]=1;ram[19][60]=0;ram[19][61]=0;ram[19][62]=1;ram[19][63]=0;ram[19][64]=0;ram[19][65]=0;ram[19][66]=1;ram[19][67]=1;ram[19][68]=1;ram[19][69]=1;ram[19][70]=1;ram[19][71]=1;ram[19][72]=1;ram[19][73]=1;ram[19][74]=1;ram[19][75]=1;ram[19][76]=1;ram[19][77]=0;ram[19][78]=1;ram[19][79]=1;ram[19][80]=1;ram[19][81]=1;ram[19][82]=1;ram[19][83]=1;ram[19][84]=1;ram[19][85]=1;ram[19][86]=0;ram[19][87]=1;ram[19][88]=1;ram[19][89]=1;ram[19][90]=1;ram[19][91]=1;ram[19][92]=1;ram[19][93]=1;ram[19][94]=1;ram[19][95]=0;ram[19][96]=1;ram[19][97]=1;ram[19][98]=0;ram[19][99]=1;ram[19][100]=1;ram[19][101]=1;ram[19][102]=1;ram[19][103]=0;ram[19][104]=1;ram[19][105]=1;ram[19][106]=1;ram[19][107]=0;ram[19][108]=1;ram[19][109]=0;ram[19][110]=0;ram[19][111]=1;ram[19][112]=1;ram[19][113]=1;ram[19][114]=1;ram[19][115]=1;ram[19][116]=0;ram[19][117]=0;ram[19][118]=1;ram[19][119]=1;ram[19][120]=0;ram[19][121]=0;ram[19][122]=1;ram[19][123]=1;ram[19][124]=1;ram[19][125]=1;ram[19][126]=1;ram[19][127]=0;ram[19][128]=1;ram[19][129]=0;ram[19][130]=1;ram[19][131]=1;ram[19][132]=0;ram[19][133]=0;ram[19][134]=1;ram[19][135]=1;ram[19][136]=0;
        ram[20][0]=1;ram[20][1]=1;ram[20][2]=1;ram[20][3]=1;ram[20][4]=1;ram[20][5]=1;ram[20][6]=1;ram[20][7]=1;ram[20][8]=0;ram[20][9]=1;ram[20][10]=1;ram[20][11]=1;ram[20][12]=1;ram[20][13]=1;ram[20][14]=0;ram[20][15]=1;ram[20][16]=1;ram[20][17]=1;ram[20][18]=1;ram[20][19]=0;ram[20][20]=1;ram[20][21]=0;ram[20][22]=0;ram[20][23]=1;ram[20][24]=1;ram[20][25]=1;ram[20][26]=1;ram[20][27]=1;ram[20][28]=0;ram[20][29]=0;ram[20][30]=1;ram[20][31]=0;ram[20][32]=1;ram[20][33]=1;ram[20][34]=1;ram[20][35]=1;ram[20][36]=1;ram[20][37]=1;ram[20][38]=0;ram[20][39]=1;ram[20][40]=1;ram[20][41]=1;ram[20][42]=0;ram[20][43]=0;ram[20][44]=1;ram[20][45]=1;ram[20][46]=0;ram[20][47]=1;ram[20][48]=0;ram[20][49]=1;ram[20][50]=0;ram[20][51]=1;ram[20][52]=0;ram[20][53]=1;ram[20][54]=1;ram[20][55]=0;ram[20][56]=0;ram[20][57]=1;ram[20][58]=1;ram[20][59]=1;ram[20][60]=0;ram[20][61]=1;ram[20][62]=1;ram[20][63]=1;ram[20][64]=0;ram[20][65]=1;ram[20][66]=1;ram[20][67]=1;ram[20][68]=1;ram[20][69]=0;ram[20][70]=1;ram[20][71]=0;ram[20][72]=1;ram[20][73]=1;ram[20][74]=0;ram[20][75]=1;ram[20][76]=1;ram[20][77]=1;ram[20][78]=0;ram[20][79]=0;ram[20][80]=0;ram[20][81]=1;ram[20][82]=1;ram[20][83]=0;ram[20][84]=0;ram[20][85]=1;ram[20][86]=0;ram[20][87]=1;ram[20][88]=1;ram[20][89]=1;ram[20][90]=0;ram[20][91]=0;ram[20][92]=0;ram[20][93]=1;ram[20][94]=0;ram[20][95]=1;ram[20][96]=1;ram[20][97]=1;ram[20][98]=1;ram[20][99]=1;ram[20][100]=1;ram[20][101]=0;ram[20][102]=1;ram[20][103]=1;ram[20][104]=0;ram[20][105]=0;ram[20][106]=1;ram[20][107]=0;ram[20][108]=1;ram[20][109]=0;ram[20][110]=1;ram[20][111]=1;ram[20][112]=1;ram[20][113]=0;ram[20][114]=0;ram[20][115]=1;ram[20][116]=1;ram[20][117]=0;ram[20][118]=1;ram[20][119]=1;ram[20][120]=1;ram[20][121]=1;ram[20][122]=0;ram[20][123]=1;ram[20][124]=0;ram[20][125]=1;ram[20][126]=0;ram[20][127]=1;ram[20][128]=1;ram[20][129]=0;ram[20][130]=0;ram[20][131]=0;ram[20][132]=1;ram[20][133]=1;ram[20][134]=1;ram[20][135]=0;ram[20][136]=1;
        ram[21][0]=1;ram[21][1]=1;ram[21][2]=1;ram[21][3]=0;ram[21][4]=1;ram[21][5]=1;ram[21][6]=1;ram[21][7]=1;ram[21][8]=0;ram[21][9]=1;ram[21][10]=0;ram[21][11]=1;ram[21][12]=0;ram[21][13]=1;ram[21][14]=0;ram[21][15]=1;ram[21][16]=1;ram[21][17]=1;ram[21][18]=1;ram[21][19]=0;ram[21][20]=0;ram[21][21]=0;ram[21][22]=1;ram[21][23]=0;ram[21][24]=1;ram[21][25]=1;ram[21][26]=0;ram[21][27]=1;ram[21][28]=1;ram[21][29]=0;ram[21][30]=0;ram[21][31]=0;ram[21][32]=0;ram[21][33]=0;ram[21][34]=1;ram[21][35]=1;ram[21][36]=0;ram[21][37]=0;ram[21][38]=1;ram[21][39]=0;ram[21][40]=0;ram[21][41]=0;ram[21][42]=0;ram[21][43]=1;ram[21][44]=1;ram[21][45]=1;ram[21][46]=1;ram[21][47]=1;ram[21][48]=0;ram[21][49]=1;ram[21][50]=1;ram[21][51]=0;ram[21][52]=0;ram[21][53]=1;ram[21][54]=1;ram[21][55]=1;ram[21][56]=1;ram[21][57]=1;ram[21][58]=0;ram[21][59]=0;ram[21][60]=1;ram[21][61]=0;ram[21][62]=0;ram[21][63]=1;ram[21][64]=0;ram[21][65]=0;ram[21][66]=1;ram[21][67]=0;ram[21][68]=1;ram[21][69]=1;ram[21][70]=1;ram[21][71]=0;ram[21][72]=1;ram[21][73]=1;ram[21][74]=0;ram[21][75]=1;ram[21][76]=0;ram[21][77]=1;ram[21][78]=1;ram[21][79]=1;ram[21][80]=1;ram[21][81]=1;ram[21][82]=1;ram[21][83]=1;ram[21][84]=0;ram[21][85]=0;ram[21][86]=0;ram[21][87]=1;ram[21][88]=1;ram[21][89]=0;ram[21][90]=1;ram[21][91]=1;ram[21][92]=1;ram[21][93]=1;ram[21][94]=0;ram[21][95]=1;ram[21][96]=1;ram[21][97]=1;ram[21][98]=0;ram[21][99]=1;ram[21][100]=1;ram[21][101]=0;ram[21][102]=0;ram[21][103]=1;ram[21][104]=1;ram[21][105]=0;ram[21][106]=1;ram[21][107]=1;ram[21][108]=1;ram[21][109]=1;ram[21][110]=0;ram[21][111]=0;ram[21][112]=1;ram[21][113]=0;ram[21][114]=1;ram[21][115]=1;ram[21][116]=1;ram[21][117]=0;ram[21][118]=1;ram[21][119]=1;ram[21][120]=1;ram[21][121]=1;ram[21][122]=1;ram[21][123]=1;ram[21][124]=1;ram[21][125]=1;ram[21][126]=1;ram[21][127]=1;ram[21][128]=1;ram[21][129]=1;ram[21][130]=1;ram[21][131]=1;ram[21][132]=0;ram[21][133]=1;ram[21][134]=1;ram[21][135]=0;ram[21][136]=1;
        ram[22][0]=1;ram[22][1]=1;ram[22][2]=1;ram[22][3]=1;ram[22][4]=1;ram[22][5]=1;ram[22][6]=1;ram[22][7]=1;ram[22][8]=1;ram[22][9]=0;ram[22][10]=1;ram[22][11]=1;ram[22][12]=1;ram[22][13]=1;ram[22][14]=0;ram[22][15]=1;ram[22][16]=1;ram[22][17]=0;ram[22][18]=1;ram[22][19]=0;ram[22][20]=1;ram[22][21]=1;ram[22][22]=1;ram[22][23]=1;ram[22][24]=1;ram[22][25]=1;ram[22][26]=0;ram[22][27]=1;ram[22][28]=1;ram[22][29]=0;ram[22][30]=0;ram[22][31]=1;ram[22][32]=1;ram[22][33]=1;ram[22][34]=0;ram[22][35]=1;ram[22][36]=1;ram[22][37]=0;ram[22][38]=1;ram[22][39]=0;ram[22][40]=1;ram[22][41]=1;ram[22][42]=1;ram[22][43]=1;ram[22][44]=1;ram[22][45]=0;ram[22][46]=1;ram[22][47]=0;ram[22][48]=1;ram[22][49]=0;ram[22][50]=0;ram[22][51]=1;ram[22][52]=1;ram[22][53]=1;ram[22][54]=1;ram[22][55]=1;ram[22][56]=0;ram[22][57]=0;ram[22][58]=1;ram[22][59]=1;ram[22][60]=1;ram[22][61]=0;ram[22][62]=1;ram[22][63]=1;ram[22][64]=1;ram[22][65]=1;ram[22][66]=0;ram[22][67]=1;ram[22][68]=1;ram[22][69]=1;ram[22][70]=1;ram[22][71]=1;ram[22][72]=1;ram[22][73]=1;ram[22][74]=1;ram[22][75]=1;ram[22][76]=0;ram[22][77]=1;ram[22][78]=0;ram[22][79]=0;ram[22][80]=0;ram[22][81]=1;ram[22][82]=1;ram[22][83]=1;ram[22][84]=1;ram[22][85]=0;ram[22][86]=0;ram[22][87]=1;ram[22][88]=1;ram[22][89]=1;ram[22][90]=1;ram[22][91]=0;ram[22][92]=0;ram[22][93]=0;ram[22][94]=1;ram[22][95]=0;ram[22][96]=1;ram[22][97]=0;ram[22][98]=0;ram[22][99]=1;ram[22][100]=0;ram[22][101]=0;ram[22][102]=0;ram[22][103]=0;ram[22][104]=1;ram[22][105]=0;ram[22][106]=0;ram[22][107]=1;ram[22][108]=0;ram[22][109]=0;ram[22][110]=1;ram[22][111]=0;ram[22][112]=0;ram[22][113]=1;ram[22][114]=1;ram[22][115]=0;ram[22][116]=1;ram[22][117]=1;ram[22][118]=1;ram[22][119]=1;ram[22][120]=1;ram[22][121]=1;ram[22][122]=1;ram[22][123]=1;ram[22][124]=0;ram[22][125]=1;ram[22][126]=1;ram[22][127]=1;ram[22][128]=1;ram[22][129]=0;ram[22][130]=0;ram[22][131]=1;ram[22][132]=1;ram[22][133]=0;ram[22][134]=1;ram[22][135]=1;ram[22][136]=0;
        ram[23][0]=1;ram[23][1]=1;ram[23][2]=0;ram[23][3]=1;ram[23][4]=0;ram[23][5]=1;ram[23][6]=0;ram[23][7]=0;ram[23][8]=1;ram[23][9]=0;ram[23][10]=1;ram[23][11]=1;ram[23][12]=1;ram[23][13]=1;ram[23][14]=1;ram[23][15]=0;ram[23][16]=0;ram[23][17]=1;ram[23][18]=1;ram[23][19]=1;ram[23][20]=1;ram[23][21]=0;ram[23][22]=0;ram[23][23]=1;ram[23][24]=0;ram[23][25]=0;ram[23][26]=1;ram[23][27]=1;ram[23][28]=1;ram[23][29]=1;ram[23][30]=1;ram[23][31]=0;ram[23][32]=1;ram[23][33]=0;ram[23][34]=1;ram[23][35]=0;ram[23][36]=1;ram[23][37]=0;ram[23][38]=1;ram[23][39]=1;ram[23][40]=0;ram[23][41]=1;ram[23][42]=0;ram[23][43]=1;ram[23][44]=0;ram[23][45]=0;ram[23][46]=1;ram[23][47]=1;ram[23][48]=0;ram[23][49]=1;ram[23][50]=1;ram[23][51]=0;ram[23][52]=1;ram[23][53]=0;ram[23][54]=1;ram[23][55]=0;ram[23][56]=1;ram[23][57]=0;ram[23][58]=0;ram[23][59]=1;ram[23][60]=0;ram[23][61]=0;ram[23][62]=0;ram[23][63]=0;ram[23][64]=1;ram[23][65]=0;ram[23][66]=0;ram[23][67]=1;ram[23][68]=1;ram[23][69]=1;ram[23][70]=1;ram[23][71]=1;ram[23][72]=1;ram[23][73]=1;ram[23][74]=0;ram[23][75]=1;ram[23][76]=1;ram[23][77]=0;ram[23][78]=1;ram[23][79]=0;ram[23][80]=1;ram[23][81]=1;ram[23][82]=1;ram[23][83]=1;ram[23][84]=1;ram[23][85]=1;ram[23][86]=1;ram[23][87]=1;ram[23][88]=1;ram[23][89]=1;ram[23][90]=1;ram[23][91]=1;ram[23][92]=0;ram[23][93]=0;ram[23][94]=1;ram[23][95]=1;ram[23][96]=1;ram[23][97]=0;ram[23][98]=1;ram[23][99]=0;ram[23][100]=1;ram[23][101]=0;ram[23][102]=1;ram[23][103]=0;ram[23][104]=1;ram[23][105]=0;ram[23][106]=0;ram[23][107]=1;ram[23][108]=0;ram[23][109]=0;ram[23][110]=0;ram[23][111]=1;ram[23][112]=0;ram[23][113]=0;ram[23][114]=0;ram[23][115]=1;ram[23][116]=1;ram[23][117]=1;ram[23][118]=1;ram[23][119]=1;ram[23][120]=0;ram[23][121]=1;ram[23][122]=1;ram[23][123]=0;ram[23][124]=0;ram[23][125]=1;ram[23][126]=1;ram[23][127]=1;ram[23][128]=0;ram[23][129]=1;ram[23][130]=0;ram[23][131]=0;ram[23][132]=1;ram[23][133]=0;ram[23][134]=1;ram[23][135]=1;ram[23][136]=0;
        ram[24][0]=0;ram[24][1]=0;ram[24][2]=1;ram[24][3]=1;ram[24][4]=0;ram[24][5]=1;ram[24][6]=1;ram[24][7]=0;ram[24][8]=1;ram[24][9]=0;ram[24][10]=0;ram[24][11]=1;ram[24][12]=1;ram[24][13]=1;ram[24][14]=1;ram[24][15]=0;ram[24][16]=1;ram[24][17]=1;ram[24][18]=1;ram[24][19]=1;ram[24][20]=1;ram[24][21]=0;ram[24][22]=0;ram[24][23]=1;ram[24][24]=1;ram[24][25]=0;ram[24][26]=1;ram[24][27]=1;ram[24][28]=1;ram[24][29]=1;ram[24][30]=0;ram[24][31]=1;ram[24][32]=0;ram[24][33]=1;ram[24][34]=1;ram[24][35]=0;ram[24][36]=1;ram[24][37]=1;ram[24][38]=1;ram[24][39]=1;ram[24][40]=0;ram[24][41]=1;ram[24][42]=1;ram[24][43]=0;ram[24][44]=1;ram[24][45]=0;ram[24][46]=1;ram[24][47]=1;ram[24][48]=0;ram[24][49]=1;ram[24][50]=1;ram[24][51]=0;ram[24][52]=0;ram[24][53]=1;ram[24][54]=1;ram[24][55]=1;ram[24][56]=1;ram[24][57]=0;ram[24][58]=1;ram[24][59]=1;ram[24][60]=1;ram[24][61]=1;ram[24][62]=0;ram[24][63]=1;ram[24][64]=1;ram[24][65]=1;ram[24][66]=0;ram[24][67]=1;ram[24][68]=0;ram[24][69]=1;ram[24][70]=1;ram[24][71]=1;ram[24][72]=1;ram[24][73]=0;ram[24][74]=1;ram[24][75]=1;ram[24][76]=1;ram[24][77]=0;ram[24][78]=1;ram[24][79]=0;ram[24][80]=0;ram[24][81]=0;ram[24][82]=1;ram[24][83]=0;ram[24][84]=0;ram[24][85]=0;ram[24][86]=0;ram[24][87]=0;ram[24][88]=1;ram[24][89]=1;ram[24][90]=0;ram[24][91]=1;ram[24][92]=0;ram[24][93]=1;ram[24][94]=1;ram[24][95]=0;ram[24][96]=0;ram[24][97]=1;ram[24][98]=0;ram[24][99]=1;ram[24][100]=0;ram[24][101]=1;ram[24][102]=1;ram[24][103]=0;ram[24][104]=0;ram[24][105]=1;ram[24][106]=1;ram[24][107]=1;ram[24][108]=0;ram[24][109]=0;ram[24][110]=1;ram[24][111]=1;ram[24][112]=1;ram[24][113]=1;ram[24][114]=1;ram[24][115]=1;ram[24][116]=0;ram[24][117]=0;ram[24][118]=1;ram[24][119]=0;ram[24][120]=1;ram[24][121]=1;ram[24][122]=1;ram[24][123]=1;ram[24][124]=1;ram[24][125]=1;ram[24][126]=0;ram[24][127]=0;ram[24][128]=0;ram[24][129]=0;ram[24][130]=1;ram[24][131]=0;ram[24][132]=0;ram[24][133]=1;ram[24][134]=1;ram[24][135]=1;ram[24][136]=0;
        ram[25][0]=1;ram[25][1]=1;ram[25][2]=1;ram[25][3]=0;ram[25][4]=0;ram[25][5]=1;ram[25][6]=1;ram[25][7]=1;ram[25][8]=1;ram[25][9]=1;ram[25][10]=0;ram[25][11]=1;ram[25][12]=0;ram[25][13]=1;ram[25][14]=1;ram[25][15]=1;ram[25][16]=0;ram[25][17]=0;ram[25][18]=1;ram[25][19]=0;ram[25][20]=0;ram[25][21]=1;ram[25][22]=1;ram[25][23]=1;ram[25][24]=1;ram[25][25]=0;ram[25][26]=1;ram[25][27]=0;ram[25][28]=1;ram[25][29]=0;ram[25][30]=1;ram[25][31]=1;ram[25][32]=1;ram[25][33]=0;ram[25][34]=1;ram[25][35]=1;ram[25][36]=0;ram[25][37]=1;ram[25][38]=0;ram[25][39]=0;ram[25][40]=0;ram[25][41]=1;ram[25][42]=0;ram[25][43]=0;ram[25][44]=0;ram[25][45]=0;ram[25][46]=1;ram[25][47]=1;ram[25][48]=1;ram[25][49]=1;ram[25][50]=1;ram[25][51]=0;ram[25][52]=1;ram[25][53]=1;ram[25][54]=0;ram[25][55]=0;ram[25][56]=1;ram[25][57]=1;ram[25][58]=1;ram[25][59]=0;ram[25][60]=1;ram[25][61]=1;ram[25][62]=0;ram[25][63]=1;ram[25][64]=1;ram[25][65]=1;ram[25][66]=0;ram[25][67]=1;ram[25][68]=1;ram[25][69]=1;ram[25][70]=0;ram[25][71]=1;ram[25][72]=1;ram[25][73]=0;ram[25][74]=0;ram[25][75]=1;ram[25][76]=0;ram[25][77]=0;ram[25][78]=0;ram[25][79]=1;ram[25][80]=1;ram[25][81]=0;ram[25][82]=0;ram[25][83]=0;ram[25][84]=0;ram[25][85]=1;ram[25][86]=0;ram[25][87]=1;ram[25][88]=1;ram[25][89]=1;ram[25][90]=1;ram[25][91]=1;ram[25][92]=1;ram[25][93]=1;ram[25][94]=0;ram[25][95]=1;ram[25][96]=1;ram[25][97]=0;ram[25][98]=0;ram[25][99]=0;ram[25][100]=1;ram[25][101]=0;ram[25][102]=0;ram[25][103]=1;ram[25][104]=0;ram[25][105]=1;ram[25][106]=0;ram[25][107]=1;ram[25][108]=1;ram[25][109]=0;ram[25][110]=0;ram[25][111]=1;ram[25][112]=1;ram[25][113]=0;ram[25][114]=0;ram[25][115]=1;ram[25][116]=1;ram[25][117]=0;ram[25][118]=1;ram[25][119]=0;ram[25][120]=0;ram[25][121]=1;ram[25][122]=1;ram[25][123]=1;ram[25][124]=1;ram[25][125]=0;ram[25][126]=1;ram[25][127]=1;ram[25][128]=1;ram[25][129]=1;ram[25][130]=0;ram[25][131]=1;ram[25][132]=1;ram[25][133]=1;ram[25][134]=1;ram[25][135]=1;ram[25][136]=0;
        ram[26][0]=0;ram[26][1]=1;ram[26][2]=0;ram[26][3]=1;ram[26][4]=1;ram[26][5]=0;ram[26][6]=1;ram[26][7]=1;ram[26][8]=1;ram[26][9]=1;ram[26][10]=0;ram[26][11]=1;ram[26][12]=0;ram[26][13]=0;ram[26][14]=1;ram[26][15]=1;ram[26][16]=1;ram[26][17]=1;ram[26][18]=0;ram[26][19]=1;ram[26][20]=1;ram[26][21]=1;ram[26][22]=1;ram[26][23]=1;ram[26][24]=1;ram[26][25]=1;ram[26][26]=0;ram[26][27]=1;ram[26][28]=1;ram[26][29]=1;ram[26][30]=1;ram[26][31]=1;ram[26][32]=1;ram[26][33]=0;ram[26][34]=1;ram[26][35]=0;ram[26][36]=1;ram[26][37]=1;ram[26][38]=1;ram[26][39]=1;ram[26][40]=1;ram[26][41]=1;ram[26][42]=1;ram[26][43]=0;ram[26][44]=1;ram[26][45]=1;ram[26][46]=1;ram[26][47]=0;ram[26][48]=1;ram[26][49]=1;ram[26][50]=1;ram[26][51]=1;ram[26][52]=1;ram[26][53]=0;ram[26][54]=1;ram[26][55]=1;ram[26][56]=1;ram[26][57]=0;ram[26][58]=1;ram[26][59]=0;ram[26][60]=1;ram[26][61]=0;ram[26][62]=0;ram[26][63]=0;ram[26][64]=0;ram[26][65]=0;ram[26][66]=1;ram[26][67]=1;ram[26][68]=1;ram[26][69]=1;ram[26][70]=0;ram[26][71]=0;ram[26][72]=0;ram[26][73]=0;ram[26][74]=1;ram[26][75]=0;ram[26][76]=0;ram[26][77]=1;ram[26][78]=0;ram[26][79]=1;ram[26][80]=1;ram[26][81]=1;ram[26][82]=0;ram[26][83]=1;ram[26][84]=1;ram[26][85]=1;ram[26][86]=1;ram[26][87]=1;ram[26][88]=1;ram[26][89]=0;ram[26][90]=0;ram[26][91]=0;ram[26][92]=1;ram[26][93]=1;ram[26][94]=1;ram[26][95]=0;ram[26][96]=0;ram[26][97]=1;ram[26][98]=1;ram[26][99]=0;ram[26][100]=1;ram[26][101]=1;ram[26][102]=0;ram[26][103]=1;ram[26][104]=1;ram[26][105]=1;ram[26][106]=0;ram[26][107]=0;ram[26][108]=0;ram[26][109]=1;ram[26][110]=1;ram[26][111]=1;ram[26][112]=1;ram[26][113]=1;ram[26][114]=1;ram[26][115]=1;ram[26][116]=1;ram[26][117]=0;ram[26][118]=1;ram[26][119]=1;ram[26][120]=1;ram[26][121]=1;ram[26][122]=1;ram[26][123]=1;ram[26][124]=0;ram[26][125]=0;ram[26][126]=0;ram[26][127]=1;ram[26][128]=1;ram[26][129]=1;ram[26][130]=0;ram[26][131]=1;ram[26][132]=1;ram[26][133]=1;ram[26][134]=1;ram[26][135]=0;ram[26][136]=0;
        ram[27][0]=1;ram[27][1]=0;ram[27][2]=0;ram[27][3]=1;ram[27][4]=1;ram[27][5]=1;ram[27][6]=0;ram[27][7]=1;ram[27][8]=1;ram[27][9]=1;ram[27][10]=0;ram[27][11]=1;ram[27][12]=0;ram[27][13]=0;ram[27][14]=0;ram[27][15]=1;ram[27][16]=1;ram[27][17]=0;ram[27][18]=0;ram[27][19]=1;ram[27][20]=0;ram[27][21]=1;ram[27][22]=0;ram[27][23]=1;ram[27][24]=1;ram[27][25]=0;ram[27][26]=1;ram[27][27]=1;ram[27][28]=1;ram[27][29]=0;ram[27][30]=1;ram[27][31]=0;ram[27][32]=0;ram[27][33]=0;ram[27][34]=0;ram[27][35]=1;ram[27][36]=0;ram[27][37]=0;ram[27][38]=0;ram[27][39]=1;ram[27][40]=0;ram[27][41]=1;ram[27][42]=1;ram[27][43]=0;ram[27][44]=1;ram[27][45]=1;ram[27][46]=1;ram[27][47]=1;ram[27][48]=0;ram[27][49]=1;ram[27][50]=1;ram[27][51]=0;ram[27][52]=1;ram[27][53]=0;ram[27][54]=0;ram[27][55]=1;ram[27][56]=0;ram[27][57]=1;ram[27][58]=1;ram[27][59]=1;ram[27][60]=0;ram[27][61]=1;ram[27][62]=0;ram[27][63]=0;ram[27][64]=1;ram[27][65]=1;ram[27][66]=1;ram[27][67]=1;ram[27][68]=0;ram[27][69]=1;ram[27][70]=1;ram[27][71]=0;ram[27][72]=1;ram[27][73]=0;ram[27][74]=1;ram[27][75]=1;ram[27][76]=1;ram[27][77]=1;ram[27][78]=1;ram[27][79]=1;ram[27][80]=1;ram[27][81]=0;ram[27][82]=0;ram[27][83]=1;ram[27][84]=1;ram[27][85]=1;ram[27][86]=1;ram[27][87]=1;ram[27][88]=1;ram[27][89]=1;ram[27][90]=1;ram[27][91]=1;ram[27][92]=1;ram[27][93]=1;ram[27][94]=0;ram[27][95]=0;ram[27][96]=0;ram[27][97]=1;ram[27][98]=1;ram[27][99]=1;ram[27][100]=0;ram[27][101]=1;ram[27][102]=0;ram[27][103]=1;ram[27][104]=1;ram[27][105]=1;ram[27][106]=0;ram[27][107]=1;ram[27][108]=1;ram[27][109]=0;ram[27][110]=0;ram[27][111]=0;ram[27][112]=1;ram[27][113]=1;ram[27][114]=1;ram[27][115]=1;ram[27][116]=1;ram[27][117]=1;ram[27][118]=1;ram[27][119]=0;ram[27][120]=0;ram[27][121]=1;ram[27][122]=1;ram[27][123]=1;ram[27][124]=0;ram[27][125]=1;ram[27][126]=1;ram[27][127]=1;ram[27][128]=1;ram[27][129]=0;ram[27][130]=0;ram[27][131]=1;ram[27][132]=1;ram[27][133]=0;ram[27][134]=0;ram[27][135]=1;ram[27][136]=1;
        ram[28][0]=1;ram[28][1]=0;ram[28][2]=0;ram[28][3]=1;ram[28][4]=0;ram[28][5]=1;ram[28][6]=1;ram[28][7]=1;ram[28][8]=1;ram[28][9]=0;ram[28][10]=1;ram[28][11]=1;ram[28][12]=1;ram[28][13]=1;ram[28][14]=0;ram[28][15]=0;ram[28][16]=1;ram[28][17]=0;ram[28][18]=0;ram[28][19]=1;ram[28][20]=1;ram[28][21]=0;ram[28][22]=0;ram[28][23]=1;ram[28][24]=0;ram[28][25]=1;ram[28][26]=1;ram[28][27]=0;ram[28][28]=1;ram[28][29]=1;ram[28][30]=1;ram[28][31]=1;ram[28][32]=1;ram[28][33]=0;ram[28][34]=1;ram[28][35]=1;ram[28][36]=0;ram[28][37]=1;ram[28][38]=0;ram[28][39]=0;ram[28][40]=1;ram[28][41]=0;ram[28][42]=0;ram[28][43]=1;ram[28][44]=1;ram[28][45]=0;ram[28][46]=1;ram[28][47]=1;ram[28][48]=1;ram[28][49]=0;ram[28][50]=0;ram[28][51]=0;ram[28][52]=1;ram[28][53]=1;ram[28][54]=1;ram[28][55]=1;ram[28][56]=1;ram[28][57]=1;ram[28][58]=1;ram[28][59]=0;ram[28][60]=1;ram[28][61]=1;ram[28][62]=0;ram[28][63]=0;ram[28][64]=0;ram[28][65]=0;ram[28][66]=1;ram[28][67]=1;ram[28][68]=1;ram[28][69]=1;ram[28][70]=1;ram[28][71]=1;ram[28][72]=0;ram[28][73]=1;ram[28][74]=1;ram[28][75]=1;ram[28][76]=0;ram[28][77]=1;ram[28][78]=1;ram[28][79]=0;ram[28][80]=1;ram[28][81]=1;ram[28][82]=0;ram[28][83]=1;ram[28][84]=1;ram[28][85]=1;ram[28][86]=1;ram[28][87]=1;ram[28][88]=1;ram[28][89]=1;ram[28][90]=1;ram[28][91]=1;ram[28][92]=1;ram[28][93]=0;ram[28][94]=0;ram[28][95]=1;ram[28][96]=1;ram[28][97]=0;ram[28][98]=1;ram[28][99]=1;ram[28][100]=1;ram[28][101]=0;ram[28][102]=1;ram[28][103]=1;ram[28][104]=1;ram[28][105]=1;ram[28][106]=0;ram[28][107]=1;ram[28][108]=1;ram[28][109]=0;ram[28][110]=1;ram[28][111]=0;ram[28][112]=1;ram[28][113]=0;ram[28][114]=0;ram[28][115]=0;ram[28][116]=1;ram[28][117]=1;ram[28][118]=0;ram[28][119]=1;ram[28][120]=1;ram[28][121]=0;ram[28][122]=1;ram[28][123]=1;ram[28][124]=1;ram[28][125]=0;ram[28][126]=0;ram[28][127]=0;ram[28][128]=1;ram[28][129]=1;ram[28][130]=1;ram[28][131]=1;ram[28][132]=1;ram[28][133]=1;ram[28][134]=0;ram[28][135]=0;ram[28][136]=1;
        ram[29][0]=1;ram[29][1]=0;ram[29][2]=1;ram[29][3]=1;ram[29][4]=1;ram[29][5]=1;ram[29][6]=0;ram[29][7]=0;ram[29][8]=0;ram[29][9]=1;ram[29][10]=1;ram[29][11]=1;ram[29][12]=0;ram[29][13]=0;ram[29][14]=0;ram[29][15]=0;ram[29][16]=1;ram[29][17]=1;ram[29][18]=0;ram[29][19]=1;ram[29][20]=1;ram[29][21]=1;ram[29][22]=0;ram[29][23]=0;ram[29][24]=0;ram[29][25]=1;ram[29][26]=1;ram[29][27]=1;ram[29][28]=1;ram[29][29]=1;ram[29][30]=1;ram[29][31]=0;ram[29][32]=1;ram[29][33]=1;ram[29][34]=1;ram[29][35]=0;ram[29][36]=1;ram[29][37]=0;ram[29][38]=1;ram[29][39]=0;ram[29][40]=1;ram[29][41]=1;ram[29][42]=0;ram[29][43]=1;ram[29][44]=1;ram[29][45]=1;ram[29][46]=1;ram[29][47]=1;ram[29][48]=1;ram[29][49]=0;ram[29][50]=1;ram[29][51]=1;ram[29][52]=1;ram[29][53]=1;ram[29][54]=1;ram[29][55]=1;ram[29][56]=0;ram[29][57]=0;ram[29][58]=1;ram[29][59]=0;ram[29][60]=0;ram[29][61]=0;ram[29][62]=0;ram[29][63]=1;ram[29][64]=1;ram[29][65]=1;ram[29][66]=1;ram[29][67]=0;ram[29][68]=1;ram[29][69]=0;ram[29][70]=0;ram[29][71]=1;ram[29][72]=0;ram[29][73]=0;ram[29][74]=1;ram[29][75]=0;ram[29][76]=0;ram[29][77]=0;ram[29][78]=1;ram[29][79]=1;ram[29][80]=0;ram[29][81]=1;ram[29][82]=1;ram[29][83]=1;ram[29][84]=1;ram[29][85]=1;ram[29][86]=1;ram[29][87]=1;ram[29][88]=0;ram[29][89]=0;ram[29][90]=1;ram[29][91]=0;ram[29][92]=1;ram[29][93]=1;ram[29][94]=1;ram[29][95]=0;ram[29][96]=1;ram[29][97]=1;ram[29][98]=1;ram[29][99]=1;ram[29][100]=1;ram[29][101]=1;ram[29][102]=1;ram[29][103]=1;ram[29][104]=1;ram[29][105]=1;ram[29][106]=1;ram[29][107]=1;ram[29][108]=1;ram[29][109]=0;ram[29][110]=1;ram[29][111]=1;ram[29][112]=1;ram[29][113]=1;ram[29][114]=1;ram[29][115]=1;ram[29][116]=1;ram[29][117]=1;ram[29][118]=1;ram[29][119]=1;ram[29][120]=0;ram[29][121]=1;ram[29][122]=1;ram[29][123]=0;ram[29][124]=1;ram[29][125]=1;ram[29][126]=1;ram[29][127]=1;ram[29][128]=1;ram[29][129]=1;ram[29][130]=0;ram[29][131]=0;ram[29][132]=0;ram[29][133]=1;ram[29][134]=1;ram[29][135]=0;ram[29][136]=1;
        ram[30][0]=0;ram[30][1]=1;ram[30][2]=0;ram[30][3]=0;ram[30][4]=1;ram[30][5]=1;ram[30][6]=1;ram[30][7]=1;ram[30][8]=0;ram[30][9]=1;ram[30][10]=0;ram[30][11]=0;ram[30][12]=0;ram[30][13]=1;ram[30][14]=0;ram[30][15]=1;ram[30][16]=1;ram[30][17]=0;ram[30][18]=1;ram[30][19]=1;ram[30][20]=1;ram[30][21]=1;ram[30][22]=1;ram[30][23]=1;ram[30][24]=0;ram[30][25]=1;ram[30][26]=1;ram[30][27]=1;ram[30][28]=1;ram[30][29]=1;ram[30][30]=1;ram[30][31]=0;ram[30][32]=1;ram[30][33]=1;ram[30][34]=1;ram[30][35]=0;ram[30][36]=1;ram[30][37]=1;ram[30][38]=1;ram[30][39]=1;ram[30][40]=1;ram[30][41]=1;ram[30][42]=0;ram[30][43]=0;ram[30][44]=1;ram[30][45]=0;ram[30][46]=1;ram[30][47]=1;ram[30][48]=1;ram[30][49]=1;ram[30][50]=1;ram[30][51]=1;ram[30][52]=1;ram[30][53]=1;ram[30][54]=0;ram[30][55]=1;ram[30][56]=0;ram[30][57]=1;ram[30][58]=1;ram[30][59]=1;ram[30][60]=1;ram[30][61]=1;ram[30][62]=0;ram[30][63]=0;ram[30][64]=1;ram[30][65]=0;ram[30][66]=1;ram[30][67]=0;ram[30][68]=0;ram[30][69]=1;ram[30][70]=0;ram[30][71]=0;ram[30][72]=1;ram[30][73]=1;ram[30][74]=0;ram[30][75]=1;ram[30][76]=1;ram[30][77]=1;ram[30][78]=1;ram[30][79]=1;ram[30][80]=0;ram[30][81]=1;ram[30][82]=0;ram[30][83]=0;ram[30][84]=1;ram[30][85]=0;ram[30][86]=0;ram[30][87]=0;ram[30][88]=0;ram[30][89]=1;ram[30][90]=1;ram[30][91]=1;ram[30][92]=1;ram[30][93]=0;ram[30][94]=0;ram[30][95]=0;ram[30][96]=0;ram[30][97]=1;ram[30][98]=1;ram[30][99]=0;ram[30][100]=1;ram[30][101]=1;ram[30][102]=1;ram[30][103]=0;ram[30][104]=1;ram[30][105]=1;ram[30][106]=1;ram[30][107]=1;ram[30][108]=1;ram[30][109]=1;ram[30][110]=1;ram[30][111]=1;ram[30][112]=1;ram[30][113]=1;ram[30][114]=1;ram[30][115]=0;ram[30][116]=1;ram[30][117]=0;ram[30][118]=0;ram[30][119]=0;ram[30][120]=1;ram[30][121]=1;ram[30][122]=1;ram[30][123]=1;ram[30][124]=0;ram[30][125]=1;ram[30][126]=0;ram[30][127]=1;ram[30][128]=1;ram[30][129]=0;ram[30][130]=0;ram[30][131]=1;ram[30][132]=1;ram[30][133]=1;ram[30][134]=1;ram[30][135]=0;ram[30][136]=0;
        ram[31][0]=1;ram[31][1]=0;ram[31][2]=1;ram[31][3]=1;ram[31][4]=1;ram[31][5]=0;ram[31][6]=1;ram[31][7]=0;ram[31][8]=0;ram[31][9]=0;ram[31][10]=0;ram[31][11]=1;ram[31][12]=1;ram[31][13]=1;ram[31][14]=1;ram[31][15]=0;ram[31][16]=0;ram[31][17]=1;ram[31][18]=0;ram[31][19]=1;ram[31][20]=1;ram[31][21]=1;ram[31][22]=0;ram[31][23]=1;ram[31][24]=1;ram[31][25]=1;ram[31][26]=1;ram[31][27]=1;ram[31][28]=1;ram[31][29]=0;ram[31][30]=1;ram[31][31]=0;ram[31][32]=1;ram[31][33]=1;ram[31][34]=1;ram[31][35]=1;ram[31][36]=1;ram[31][37]=1;ram[31][38]=1;ram[31][39]=1;ram[31][40]=1;ram[31][41]=1;ram[31][42]=1;ram[31][43]=1;ram[31][44]=1;ram[31][45]=1;ram[31][46]=1;ram[31][47]=1;ram[31][48]=1;ram[31][49]=1;ram[31][50]=1;ram[31][51]=1;ram[31][52]=0;ram[31][53]=0;ram[31][54]=0;ram[31][55]=1;ram[31][56]=0;ram[31][57]=0;ram[31][58]=1;ram[31][59]=0;ram[31][60]=1;ram[31][61]=1;ram[31][62]=0;ram[31][63]=1;ram[31][64]=1;ram[31][65]=1;ram[31][66]=1;ram[31][67]=1;ram[31][68]=1;ram[31][69]=1;ram[31][70]=0;ram[31][71]=1;ram[31][72]=1;ram[31][73]=1;ram[31][74]=1;ram[31][75]=1;ram[31][76]=0;ram[31][77]=0;ram[31][78]=1;ram[31][79]=1;ram[31][80]=0;ram[31][81]=0;ram[31][82]=1;ram[31][83]=1;ram[31][84]=1;ram[31][85]=1;ram[31][86]=1;ram[31][87]=0;ram[31][88]=0;ram[31][89]=0;ram[31][90]=1;ram[31][91]=1;ram[31][92]=0;ram[31][93]=1;ram[31][94]=1;ram[31][95]=0;ram[31][96]=1;ram[31][97]=1;ram[31][98]=1;ram[31][99]=0;ram[31][100]=1;ram[31][101]=1;ram[31][102]=1;ram[31][103]=0;ram[31][104]=1;ram[31][105]=0;ram[31][106]=1;ram[31][107]=0;ram[31][108]=0;ram[31][109]=0;ram[31][110]=1;ram[31][111]=0;ram[31][112]=0;ram[31][113]=1;ram[31][114]=1;ram[31][115]=1;ram[31][116]=1;ram[31][117]=1;ram[31][118]=0;ram[31][119]=1;ram[31][120]=1;ram[31][121]=1;ram[31][122]=0;ram[31][123]=0;ram[31][124]=1;ram[31][125]=1;ram[31][126]=1;ram[31][127]=0;ram[31][128]=1;ram[31][129]=1;ram[31][130]=1;ram[31][131]=0;ram[31][132]=1;ram[31][133]=1;ram[31][134]=1;ram[31][135]=1;ram[31][136]=0;
        ram[32][0]=1;ram[32][1]=1;ram[32][2]=0;ram[32][3]=0;ram[32][4]=1;ram[32][5]=0;ram[32][6]=1;ram[32][7]=0;ram[32][8]=0;ram[32][9]=0;ram[32][10]=0;ram[32][11]=0;ram[32][12]=0;ram[32][13]=1;ram[32][14]=1;ram[32][15]=1;ram[32][16]=0;ram[32][17]=1;ram[32][18]=1;ram[32][19]=1;ram[32][20]=1;ram[32][21]=0;ram[32][22]=0;ram[32][23]=1;ram[32][24]=1;ram[32][25]=0;ram[32][26]=1;ram[32][27]=1;ram[32][28]=0;ram[32][29]=0;ram[32][30]=1;ram[32][31]=1;ram[32][32]=0;ram[32][33]=1;ram[32][34]=1;ram[32][35]=1;ram[32][36]=0;ram[32][37]=0;ram[32][38]=0;ram[32][39]=1;ram[32][40]=1;ram[32][41]=1;ram[32][42]=1;ram[32][43]=1;ram[32][44]=0;ram[32][45]=1;ram[32][46]=1;ram[32][47]=0;ram[32][48]=0;ram[32][49]=1;ram[32][50]=0;ram[32][51]=0;ram[32][52]=1;ram[32][53]=1;ram[32][54]=0;ram[32][55]=1;ram[32][56]=1;ram[32][57]=1;ram[32][58]=1;ram[32][59]=1;ram[32][60]=1;ram[32][61]=1;ram[32][62]=1;ram[32][63]=1;ram[32][64]=1;ram[32][65]=1;ram[32][66]=0;ram[32][67]=1;ram[32][68]=1;ram[32][69]=1;ram[32][70]=1;ram[32][71]=1;ram[32][72]=1;ram[32][73]=0;ram[32][74]=0;ram[32][75]=1;ram[32][76]=0;ram[32][77]=1;ram[32][78]=1;ram[32][79]=0;ram[32][80]=1;ram[32][81]=1;ram[32][82]=1;ram[32][83]=1;ram[32][84]=1;ram[32][85]=1;ram[32][86]=1;ram[32][87]=1;ram[32][88]=1;ram[32][89]=1;ram[32][90]=0;ram[32][91]=0;ram[32][92]=0;ram[32][93]=0;ram[32][94]=0;ram[32][95]=1;ram[32][96]=1;ram[32][97]=1;ram[32][98]=0;ram[32][99]=1;ram[32][100]=0;ram[32][101]=1;ram[32][102]=1;ram[32][103]=1;ram[32][104]=1;ram[32][105]=1;ram[32][106]=1;ram[32][107]=1;ram[32][108]=1;ram[32][109]=1;ram[32][110]=1;ram[32][111]=1;ram[32][112]=1;ram[32][113]=1;ram[32][114]=0;ram[32][115]=1;ram[32][116]=1;ram[32][117]=1;ram[32][118]=0;ram[32][119]=1;ram[32][120]=1;ram[32][121]=1;ram[32][122]=0;ram[32][123]=1;ram[32][124]=1;ram[32][125]=1;ram[32][126]=1;ram[32][127]=1;ram[32][128]=1;ram[32][129]=0;ram[32][130]=0;ram[32][131]=1;ram[32][132]=1;ram[32][133]=0;ram[32][134]=1;ram[32][135]=0;ram[32][136]=1;
        ram[33][0]=0;ram[33][1]=1;ram[33][2]=0;ram[33][3]=1;ram[33][4]=1;ram[33][5]=1;ram[33][6]=0;ram[33][7]=0;ram[33][8]=1;ram[33][9]=0;ram[33][10]=0;ram[33][11]=0;ram[33][12]=0;ram[33][13]=1;ram[33][14]=1;ram[33][15]=1;ram[33][16]=1;ram[33][17]=0;ram[33][18]=0;ram[33][19]=1;ram[33][20]=1;ram[33][21]=0;ram[33][22]=1;ram[33][23]=1;ram[33][24]=1;ram[33][25]=0;ram[33][26]=1;ram[33][27]=1;ram[33][28]=1;ram[33][29]=1;ram[33][30]=1;ram[33][31]=1;ram[33][32]=1;ram[33][33]=1;ram[33][34]=1;ram[33][35]=1;ram[33][36]=1;ram[33][37]=1;ram[33][38]=0;ram[33][39]=0;ram[33][40]=1;ram[33][41]=1;ram[33][42]=0;ram[33][43]=0;ram[33][44]=1;ram[33][45]=1;ram[33][46]=0;ram[33][47]=1;ram[33][48]=1;ram[33][49]=1;ram[33][50]=1;ram[33][51]=1;ram[33][52]=1;ram[33][53]=0;ram[33][54]=1;ram[33][55]=0;ram[33][56]=1;ram[33][57]=0;ram[33][58]=1;ram[33][59]=1;ram[33][60]=1;ram[33][61]=0;ram[33][62]=0;ram[33][63]=1;ram[33][64]=1;ram[33][65]=1;ram[33][66]=0;ram[33][67]=1;ram[33][68]=1;ram[33][69]=1;ram[33][70]=1;ram[33][71]=1;ram[33][72]=1;ram[33][73]=0;ram[33][74]=1;ram[33][75]=1;ram[33][76]=1;ram[33][77]=1;ram[33][78]=0;ram[33][79]=0;ram[33][80]=0;ram[33][81]=1;ram[33][82]=1;ram[33][83]=1;ram[33][84]=1;ram[33][85]=1;ram[33][86]=0;ram[33][87]=1;ram[33][88]=0;ram[33][89]=1;ram[33][90]=1;ram[33][91]=1;ram[33][92]=1;ram[33][93]=0;ram[33][94]=0;ram[33][95]=1;ram[33][96]=1;ram[33][97]=1;ram[33][98]=1;ram[33][99]=1;ram[33][100]=1;ram[33][101]=0;ram[33][102]=1;ram[33][103]=0;ram[33][104]=0;ram[33][105]=1;ram[33][106]=1;ram[33][107]=1;ram[33][108]=1;ram[33][109]=1;ram[33][110]=0;ram[33][111]=1;ram[33][112]=1;ram[33][113]=1;ram[33][114]=1;ram[33][115]=1;ram[33][116]=0;ram[33][117]=0;ram[33][118]=1;ram[33][119]=1;ram[33][120]=1;ram[33][121]=1;ram[33][122]=1;ram[33][123]=1;ram[33][124]=0;ram[33][125]=1;ram[33][126]=0;ram[33][127]=1;ram[33][128]=1;ram[33][129]=1;ram[33][130]=1;ram[33][131]=1;ram[33][132]=1;ram[33][133]=1;ram[33][134]=1;ram[33][135]=1;ram[33][136]=0;
        ram[34][0]=1;ram[34][1]=0;ram[34][2]=0;ram[34][3]=1;ram[34][4]=1;ram[34][5]=1;ram[34][6]=1;ram[34][7]=0;ram[34][8]=1;ram[34][9]=1;ram[34][10]=1;ram[34][11]=1;ram[34][12]=0;ram[34][13]=1;ram[34][14]=0;ram[34][15]=1;ram[34][16]=0;ram[34][17]=1;ram[34][18]=1;ram[34][19]=0;ram[34][20]=0;ram[34][21]=1;ram[34][22]=1;ram[34][23]=0;ram[34][24]=1;ram[34][25]=1;ram[34][26]=1;ram[34][27]=1;ram[34][28]=1;ram[34][29]=1;ram[34][30]=1;ram[34][31]=1;ram[34][32]=1;ram[34][33]=1;ram[34][34]=1;ram[34][35]=0;ram[34][36]=1;ram[34][37]=0;ram[34][38]=0;ram[34][39]=0;ram[34][40]=1;ram[34][41]=0;ram[34][42]=1;ram[34][43]=0;ram[34][44]=1;ram[34][45]=0;ram[34][46]=1;ram[34][47]=0;ram[34][48]=1;ram[34][49]=0;ram[34][50]=1;ram[34][51]=1;ram[34][52]=1;ram[34][53]=1;ram[34][54]=1;ram[34][55]=1;ram[34][56]=1;ram[34][57]=0;ram[34][58]=1;ram[34][59]=0;ram[34][60]=1;ram[34][61]=1;ram[34][62]=0;ram[34][63]=0;ram[34][64]=0;ram[34][65]=1;ram[34][66]=1;ram[34][67]=1;ram[34][68]=1;ram[34][69]=0;ram[34][70]=0;ram[34][71]=0;ram[34][72]=1;ram[34][73]=0;ram[34][74]=1;ram[34][75]=1;ram[34][76]=1;ram[34][77]=1;ram[34][78]=0;ram[34][79]=0;ram[34][80]=0;ram[34][81]=1;ram[34][82]=1;ram[34][83]=0;ram[34][84]=1;ram[34][85]=1;ram[34][86]=0;ram[34][87]=0;ram[34][88]=1;ram[34][89]=1;ram[34][90]=1;ram[34][91]=0;ram[34][92]=1;ram[34][93]=1;ram[34][94]=1;ram[34][95]=0;ram[34][96]=1;ram[34][97]=1;ram[34][98]=0;ram[34][99]=1;ram[34][100]=0;ram[34][101]=1;ram[34][102]=0;ram[34][103]=1;ram[34][104]=1;ram[34][105]=1;ram[34][106]=1;ram[34][107]=1;ram[34][108]=1;ram[34][109]=1;ram[34][110]=1;ram[34][111]=0;ram[34][112]=1;ram[34][113]=1;ram[34][114]=1;ram[34][115]=1;ram[34][116]=0;ram[34][117]=1;ram[34][118]=1;ram[34][119]=0;ram[34][120]=0;ram[34][121]=0;ram[34][122]=1;ram[34][123]=1;ram[34][124]=1;ram[34][125]=1;ram[34][126]=1;ram[34][127]=1;ram[34][128]=0;ram[34][129]=0;ram[34][130]=1;ram[34][131]=1;ram[34][132]=1;ram[34][133]=0;ram[34][134]=0;ram[34][135]=1;ram[34][136]=1;
        ram[35][0]=0;ram[35][1]=1;ram[35][2]=1;ram[35][3]=1;ram[35][4]=1;ram[35][5]=1;ram[35][6]=0;ram[35][7]=1;ram[35][8]=0;ram[35][9]=1;ram[35][10]=1;ram[35][11]=1;ram[35][12]=0;ram[35][13]=1;ram[35][14]=1;ram[35][15]=1;ram[35][16]=1;ram[35][17]=0;ram[35][18]=1;ram[35][19]=1;ram[35][20]=1;ram[35][21]=1;ram[35][22]=1;ram[35][23]=1;ram[35][24]=1;ram[35][25]=1;ram[35][26]=1;ram[35][27]=1;ram[35][28]=1;ram[35][29]=1;ram[35][30]=0;ram[35][31]=1;ram[35][32]=1;ram[35][33]=0;ram[35][34]=1;ram[35][35]=1;ram[35][36]=1;ram[35][37]=0;ram[35][38]=1;ram[35][39]=1;ram[35][40]=0;ram[35][41]=0;ram[35][42]=1;ram[35][43]=0;ram[35][44]=0;ram[35][45]=1;ram[35][46]=1;ram[35][47]=1;ram[35][48]=1;ram[35][49]=1;ram[35][50]=1;ram[35][51]=0;ram[35][52]=0;ram[35][53]=1;ram[35][54]=0;ram[35][55]=0;ram[35][56]=1;ram[35][57]=1;ram[35][58]=0;ram[35][59]=0;ram[35][60]=1;ram[35][61]=1;ram[35][62]=1;ram[35][63]=1;ram[35][64]=0;ram[35][65]=0;ram[35][66]=1;ram[35][67]=1;ram[35][68]=1;ram[35][69]=1;ram[35][70]=0;ram[35][71]=1;ram[35][72]=1;ram[35][73]=0;ram[35][74]=0;ram[35][75]=1;ram[35][76]=1;ram[35][77]=1;ram[35][78]=1;ram[35][79]=1;ram[35][80]=1;ram[35][81]=0;ram[35][82]=0;ram[35][83]=1;ram[35][84]=1;ram[35][85]=1;ram[35][86]=1;ram[35][87]=1;ram[35][88]=1;ram[35][89]=0;ram[35][90]=1;ram[35][91]=1;ram[35][92]=0;ram[35][93]=1;ram[35][94]=1;ram[35][95]=1;ram[35][96]=0;ram[35][97]=1;ram[35][98]=1;ram[35][99]=1;ram[35][100]=1;ram[35][101]=1;ram[35][102]=1;ram[35][103]=1;ram[35][104]=1;ram[35][105]=0;ram[35][106]=0;ram[35][107]=1;ram[35][108]=0;ram[35][109]=0;ram[35][110]=1;ram[35][111]=1;ram[35][112]=0;ram[35][113]=1;ram[35][114]=1;ram[35][115]=0;ram[35][116]=1;ram[35][117]=1;ram[35][118]=1;ram[35][119]=0;ram[35][120]=1;ram[35][121]=1;ram[35][122]=1;ram[35][123]=1;ram[35][124]=1;ram[35][125]=1;ram[35][126]=1;ram[35][127]=1;ram[35][128]=1;ram[35][129]=1;ram[35][130]=0;ram[35][131]=0;ram[35][132]=0;ram[35][133]=0;ram[35][134]=1;ram[35][135]=1;ram[35][136]=0;
        ram[36][0]=1;ram[36][1]=1;ram[36][2]=1;ram[36][3]=0;ram[36][4]=1;ram[36][5]=1;ram[36][6]=1;ram[36][7]=0;ram[36][8]=1;ram[36][9]=1;ram[36][10]=1;ram[36][11]=1;ram[36][12]=1;ram[36][13]=1;ram[36][14]=1;ram[36][15]=1;ram[36][16]=1;ram[36][17]=1;ram[36][18]=0;ram[36][19]=0;ram[36][20]=0;ram[36][21]=1;ram[36][22]=0;ram[36][23]=1;ram[36][24]=0;ram[36][25]=0;ram[36][26]=1;ram[36][27]=1;ram[36][28]=1;ram[36][29]=0;ram[36][30]=1;ram[36][31]=0;ram[36][32]=1;ram[36][33]=1;ram[36][34]=0;ram[36][35]=1;ram[36][36]=1;ram[36][37]=0;ram[36][38]=1;ram[36][39]=1;ram[36][40]=1;ram[36][41]=1;ram[36][42]=1;ram[36][43]=0;ram[36][44]=0;ram[36][45]=1;ram[36][46]=1;ram[36][47]=1;ram[36][48]=1;ram[36][49]=1;ram[36][50]=0;ram[36][51]=1;ram[36][52]=1;ram[36][53]=1;ram[36][54]=1;ram[36][55]=0;ram[36][56]=1;ram[36][57]=0;ram[36][58]=1;ram[36][59]=1;ram[36][60]=0;ram[36][61]=1;ram[36][62]=0;ram[36][63]=1;ram[36][64]=1;ram[36][65]=1;ram[36][66]=1;ram[36][67]=0;ram[36][68]=0;ram[36][69]=1;ram[36][70]=1;ram[36][71]=1;ram[36][72]=0;ram[36][73]=0;ram[36][74]=1;ram[36][75]=0;ram[36][76]=1;ram[36][77]=0;ram[36][78]=0;ram[36][79]=1;ram[36][80]=0;ram[36][81]=1;ram[36][82]=1;ram[36][83]=1;ram[36][84]=1;ram[36][85]=1;ram[36][86]=1;ram[36][87]=0;ram[36][88]=1;ram[36][89]=0;ram[36][90]=1;ram[36][91]=1;ram[36][92]=1;ram[36][93]=1;ram[36][94]=1;ram[36][95]=1;ram[36][96]=0;ram[36][97]=1;ram[36][98]=0;ram[36][99]=1;ram[36][100]=0;ram[36][101]=1;ram[36][102]=0;ram[36][103]=1;ram[36][104]=1;ram[36][105]=1;ram[36][106]=1;ram[36][107]=1;ram[36][108]=0;ram[36][109]=0;ram[36][110]=0;ram[36][111]=1;ram[36][112]=1;ram[36][113]=0;ram[36][114]=1;ram[36][115]=1;ram[36][116]=1;ram[36][117]=1;ram[36][118]=1;ram[36][119]=0;ram[36][120]=1;ram[36][121]=1;ram[36][122]=1;ram[36][123]=1;ram[36][124]=1;ram[36][125]=1;ram[36][126]=1;ram[36][127]=1;ram[36][128]=1;ram[36][129]=1;ram[36][130]=1;ram[36][131]=1;ram[36][132]=1;ram[36][133]=1;ram[36][134]=1;ram[36][135]=1;ram[36][136]=1;
        ram[37][0]=1;ram[37][1]=1;ram[37][2]=1;ram[37][3]=0;ram[37][4]=1;ram[37][5]=1;ram[37][6]=0;ram[37][7]=1;ram[37][8]=1;ram[37][9]=1;ram[37][10]=0;ram[37][11]=0;ram[37][12]=0;ram[37][13]=1;ram[37][14]=0;ram[37][15]=0;ram[37][16]=1;ram[37][17]=0;ram[37][18]=0;ram[37][19]=1;ram[37][20]=0;ram[37][21]=1;ram[37][22]=1;ram[37][23]=1;ram[37][24]=0;ram[37][25]=1;ram[37][26]=1;ram[37][27]=1;ram[37][28]=1;ram[37][29]=0;ram[37][30]=1;ram[37][31]=0;ram[37][32]=1;ram[37][33]=1;ram[37][34]=1;ram[37][35]=1;ram[37][36]=0;ram[37][37]=0;ram[37][38]=1;ram[37][39]=1;ram[37][40]=1;ram[37][41]=0;ram[37][42]=0;ram[37][43]=1;ram[37][44]=1;ram[37][45]=0;ram[37][46]=1;ram[37][47]=1;ram[37][48]=1;ram[37][49]=1;ram[37][50]=1;ram[37][51]=1;ram[37][52]=0;ram[37][53]=1;ram[37][54]=1;ram[37][55]=1;ram[37][56]=1;ram[37][57]=1;ram[37][58]=1;ram[37][59]=1;ram[37][60]=1;ram[37][61]=0;ram[37][62]=1;ram[37][63]=1;ram[37][64]=1;ram[37][65]=1;ram[37][66]=1;ram[37][67]=1;ram[37][68]=1;ram[37][69]=1;ram[37][70]=1;ram[37][71]=1;ram[37][72]=1;ram[37][73]=1;ram[37][74]=1;ram[37][75]=0;ram[37][76]=0;ram[37][77]=0;ram[37][78]=1;ram[37][79]=0;ram[37][80]=1;ram[37][81]=0;ram[37][82]=0;ram[37][83]=0;ram[37][84]=1;ram[37][85]=0;ram[37][86]=1;ram[37][87]=0;ram[37][88]=1;ram[37][89]=0;ram[37][90]=1;ram[37][91]=1;ram[37][92]=1;ram[37][93]=1;ram[37][94]=1;ram[37][95]=1;ram[37][96]=1;ram[37][97]=1;ram[37][98]=0;ram[37][99]=1;ram[37][100]=1;ram[37][101]=0;ram[37][102]=1;ram[37][103]=0;ram[37][104]=0;ram[37][105]=1;ram[37][106]=1;ram[37][107]=0;ram[37][108]=1;ram[37][109]=0;ram[37][110]=0;ram[37][111]=1;ram[37][112]=1;ram[37][113]=1;ram[37][114]=1;ram[37][115]=0;ram[37][116]=0;ram[37][117]=1;ram[37][118]=1;ram[37][119]=1;ram[37][120]=1;ram[37][121]=1;ram[37][122]=1;ram[37][123]=0;ram[37][124]=1;ram[37][125]=1;ram[37][126]=1;ram[37][127]=1;ram[37][128]=1;ram[37][129]=1;ram[37][130]=1;ram[37][131]=1;ram[37][132]=1;ram[37][133]=1;ram[37][134]=1;ram[37][135]=0;ram[37][136]=1;
        ram[38][0]=0;ram[38][1]=1;ram[38][2]=0;ram[38][3]=0;ram[38][4]=1;ram[38][5]=0;ram[38][6]=1;ram[38][7]=0;ram[38][8]=1;ram[38][9]=1;ram[38][10]=1;ram[38][11]=1;ram[38][12]=1;ram[38][13]=0;ram[38][14]=1;ram[38][15]=1;ram[38][16]=1;ram[38][17]=0;ram[38][18]=1;ram[38][19]=0;ram[38][20]=1;ram[38][21]=1;ram[38][22]=1;ram[38][23]=0;ram[38][24]=0;ram[38][25]=1;ram[38][26]=1;ram[38][27]=1;ram[38][28]=1;ram[38][29]=1;ram[38][30]=0;ram[38][31]=1;ram[38][32]=0;ram[38][33]=0;ram[38][34]=1;ram[38][35]=1;ram[38][36]=1;ram[38][37]=1;ram[38][38]=1;ram[38][39]=1;ram[38][40]=1;ram[38][41]=1;ram[38][42]=1;ram[38][43]=1;ram[38][44]=0;ram[38][45]=0;ram[38][46]=1;ram[38][47]=0;ram[38][48]=1;ram[38][49]=1;ram[38][50]=1;ram[38][51]=1;ram[38][52]=1;ram[38][53]=0;ram[38][54]=0;ram[38][55]=0;ram[38][56]=1;ram[38][57]=1;ram[38][58]=1;ram[38][59]=1;ram[38][60]=1;ram[38][61]=1;ram[38][62]=1;ram[38][63]=1;ram[38][64]=1;ram[38][65]=1;ram[38][66]=0;ram[38][67]=0;ram[38][68]=1;ram[38][69]=0;ram[38][70]=0;ram[38][71]=1;ram[38][72]=1;ram[38][73]=1;ram[38][74]=0;ram[38][75]=0;ram[38][76]=0;ram[38][77]=1;ram[38][78]=1;ram[38][79]=1;ram[38][80]=1;ram[38][81]=1;ram[38][82]=0;ram[38][83]=1;ram[38][84]=1;ram[38][85]=1;ram[38][86]=0;ram[38][87]=0;ram[38][88]=1;ram[38][89]=1;ram[38][90]=1;ram[38][91]=1;ram[38][92]=1;ram[38][93]=1;ram[38][94]=1;ram[38][95]=0;ram[38][96]=1;ram[38][97]=0;ram[38][98]=1;ram[38][99]=0;ram[38][100]=0;ram[38][101]=0;ram[38][102]=1;ram[38][103]=1;ram[38][104]=1;ram[38][105]=0;ram[38][106]=0;ram[38][107]=1;ram[38][108]=0;ram[38][109]=1;ram[38][110]=0;ram[38][111]=0;ram[38][112]=0;ram[38][113]=1;ram[38][114]=0;ram[38][115]=1;ram[38][116]=1;ram[38][117]=0;ram[38][118]=1;ram[38][119]=1;ram[38][120]=1;ram[38][121]=1;ram[38][122]=0;ram[38][123]=1;ram[38][124]=1;ram[38][125]=1;ram[38][126]=1;ram[38][127]=1;ram[38][128]=0;ram[38][129]=0;ram[38][130]=1;ram[38][131]=1;ram[38][132]=0;ram[38][133]=1;ram[38][134]=0;ram[38][135]=1;ram[38][136]=1;
        ram[39][0]=1;ram[39][1]=0;ram[39][2]=0;ram[39][3]=1;ram[39][4]=1;ram[39][5]=1;ram[39][6]=0;ram[39][7]=1;ram[39][8]=1;ram[39][9]=1;ram[39][10]=1;ram[39][11]=1;ram[39][12]=1;ram[39][13]=0;ram[39][14]=1;ram[39][15]=1;ram[39][16]=1;ram[39][17]=0;ram[39][18]=1;ram[39][19]=1;ram[39][20]=1;ram[39][21]=1;ram[39][22]=1;ram[39][23]=1;ram[39][24]=1;ram[39][25]=1;ram[39][26]=1;ram[39][27]=1;ram[39][28]=0;ram[39][29]=1;ram[39][30]=1;ram[39][31]=1;ram[39][32]=0;ram[39][33]=1;ram[39][34]=1;ram[39][35]=1;ram[39][36]=1;ram[39][37]=1;ram[39][38]=1;ram[39][39]=0;ram[39][40]=1;ram[39][41]=1;ram[39][42]=1;ram[39][43]=1;ram[39][44]=1;ram[39][45]=0;ram[39][46]=0;ram[39][47]=1;ram[39][48]=1;ram[39][49]=1;ram[39][50]=1;ram[39][51]=1;ram[39][52]=1;ram[39][53]=1;ram[39][54]=1;ram[39][55]=1;ram[39][56]=0;ram[39][57]=1;ram[39][58]=1;ram[39][59]=0;ram[39][60]=1;ram[39][61]=0;ram[39][62]=0;ram[39][63]=1;ram[39][64]=1;ram[39][65]=0;ram[39][66]=1;ram[39][67]=1;ram[39][68]=1;ram[39][69]=1;ram[39][70]=1;ram[39][71]=0;ram[39][72]=1;ram[39][73]=1;ram[39][74]=0;ram[39][75]=0;ram[39][76]=0;ram[39][77]=1;ram[39][78]=1;ram[39][79]=0;ram[39][80]=1;ram[39][81]=1;ram[39][82]=1;ram[39][83]=1;ram[39][84]=1;ram[39][85]=1;ram[39][86]=0;ram[39][87]=1;ram[39][88]=1;ram[39][89]=1;ram[39][90]=1;ram[39][91]=1;ram[39][92]=1;ram[39][93]=0;ram[39][94]=0;ram[39][95]=1;ram[39][96]=1;ram[39][97]=1;ram[39][98]=1;ram[39][99]=0;ram[39][100]=1;ram[39][101]=1;ram[39][102]=1;ram[39][103]=1;ram[39][104]=1;ram[39][105]=1;ram[39][106]=1;ram[39][107]=0;ram[39][108]=1;ram[39][109]=1;ram[39][110]=1;ram[39][111]=1;ram[39][112]=1;ram[39][113]=0;ram[39][114]=0;ram[39][115]=1;ram[39][116]=1;ram[39][117]=1;ram[39][118]=0;ram[39][119]=1;ram[39][120]=1;ram[39][121]=1;ram[39][122]=1;ram[39][123]=0;ram[39][124]=1;ram[39][125]=1;ram[39][126]=0;ram[39][127]=1;ram[39][128]=1;ram[39][129]=1;ram[39][130]=1;ram[39][131]=0;ram[39][132]=1;ram[39][133]=1;ram[39][134]=0;ram[39][135]=1;ram[39][136]=0;
        ram[40][0]=1;ram[40][1]=0;ram[40][2]=1;ram[40][3]=1;ram[40][4]=0;ram[40][5]=1;ram[40][6]=1;ram[40][7]=1;ram[40][8]=0;ram[40][9]=1;ram[40][10]=0;ram[40][11]=1;ram[40][12]=0;ram[40][13]=0;ram[40][14]=1;ram[40][15]=0;ram[40][16]=1;ram[40][17]=1;ram[40][18]=0;ram[40][19]=0;ram[40][20]=1;ram[40][21]=0;ram[40][22]=1;ram[40][23]=1;ram[40][24]=0;ram[40][25]=0;ram[40][26]=1;ram[40][27]=1;ram[40][28]=1;ram[40][29]=1;ram[40][30]=1;ram[40][31]=0;ram[40][32]=1;ram[40][33]=1;ram[40][34]=1;ram[40][35]=1;ram[40][36]=0;ram[40][37]=1;ram[40][38]=0;ram[40][39]=1;ram[40][40]=0;ram[40][41]=0;ram[40][42]=1;ram[40][43]=0;ram[40][44]=1;ram[40][45]=1;ram[40][46]=0;ram[40][47]=1;ram[40][48]=0;ram[40][49]=1;ram[40][50]=1;ram[40][51]=1;ram[40][52]=1;ram[40][53]=1;ram[40][54]=0;ram[40][55]=0;ram[40][56]=1;ram[40][57]=1;ram[40][58]=0;ram[40][59]=1;ram[40][60]=0;ram[40][61]=1;ram[40][62]=1;ram[40][63]=1;ram[40][64]=1;ram[40][65]=1;ram[40][66]=0;ram[40][67]=1;ram[40][68]=1;ram[40][69]=1;ram[40][70]=0;ram[40][71]=1;ram[40][72]=1;ram[40][73]=0;ram[40][74]=1;ram[40][75]=1;ram[40][76]=1;ram[40][77]=1;ram[40][78]=0;ram[40][79]=0;ram[40][80]=1;ram[40][81]=1;ram[40][82]=0;ram[40][83]=0;ram[40][84]=1;ram[40][85]=0;ram[40][86]=0;ram[40][87]=1;ram[40][88]=0;ram[40][89]=1;ram[40][90]=0;ram[40][91]=0;ram[40][92]=0;ram[40][93]=1;ram[40][94]=1;ram[40][95]=0;ram[40][96]=0;ram[40][97]=1;ram[40][98]=1;ram[40][99]=1;ram[40][100]=0;ram[40][101]=1;ram[40][102]=1;ram[40][103]=1;ram[40][104]=0;ram[40][105]=1;ram[40][106]=1;ram[40][107]=1;ram[40][108]=1;ram[40][109]=0;ram[40][110]=0;ram[40][111]=1;ram[40][112]=0;ram[40][113]=1;ram[40][114]=1;ram[40][115]=1;ram[40][116]=0;ram[40][117]=1;ram[40][118]=1;ram[40][119]=0;ram[40][120]=1;ram[40][121]=0;ram[40][122]=0;ram[40][123]=1;ram[40][124]=1;ram[40][125]=1;ram[40][126]=1;ram[40][127]=1;ram[40][128]=1;ram[40][129]=1;ram[40][130]=1;ram[40][131]=1;ram[40][132]=1;ram[40][133]=0;ram[40][134]=1;ram[40][135]=0;ram[40][136]=0;
        ram[41][0]=1;ram[41][1]=1;ram[41][2]=0;ram[41][3]=1;ram[41][4]=0;ram[41][5]=1;ram[41][6]=1;ram[41][7]=0;ram[41][8]=1;ram[41][9]=0;ram[41][10]=1;ram[41][11]=1;ram[41][12]=0;ram[41][13]=1;ram[41][14]=1;ram[41][15]=0;ram[41][16]=1;ram[41][17]=0;ram[41][18]=1;ram[41][19]=1;ram[41][20]=1;ram[41][21]=1;ram[41][22]=1;ram[41][23]=1;ram[41][24]=1;ram[41][25]=1;ram[41][26]=1;ram[41][27]=1;ram[41][28]=1;ram[41][29]=0;ram[41][30]=0;ram[41][31]=1;ram[41][32]=0;ram[41][33]=0;ram[41][34]=1;ram[41][35]=1;ram[41][36]=0;ram[41][37]=1;ram[41][38]=1;ram[41][39]=0;ram[41][40]=1;ram[41][41]=0;ram[41][42]=0;ram[41][43]=1;ram[41][44]=1;ram[41][45]=0;ram[41][46]=1;ram[41][47]=1;ram[41][48]=1;ram[41][49]=1;ram[41][50]=0;ram[41][51]=1;ram[41][52]=0;ram[41][53]=1;ram[41][54]=0;ram[41][55]=1;ram[41][56]=1;ram[41][57]=1;ram[41][58]=1;ram[41][59]=1;ram[41][60]=1;ram[41][61]=0;ram[41][62]=1;ram[41][63]=0;ram[41][64]=1;ram[41][65]=1;ram[41][66]=1;ram[41][67]=1;ram[41][68]=1;ram[41][69]=1;ram[41][70]=1;ram[41][71]=1;ram[41][72]=1;ram[41][73]=1;ram[41][74]=1;ram[41][75]=1;ram[41][76]=1;ram[41][77]=1;ram[41][78]=1;ram[41][79]=1;ram[41][80]=0;ram[41][81]=0;ram[41][82]=1;ram[41][83]=1;ram[41][84]=0;ram[41][85]=0;ram[41][86]=1;ram[41][87]=1;ram[41][88]=0;ram[41][89]=1;ram[41][90]=0;ram[41][91]=1;ram[41][92]=1;ram[41][93]=1;ram[41][94]=1;ram[41][95]=1;ram[41][96]=0;ram[41][97]=1;ram[41][98]=0;ram[41][99]=0;ram[41][100]=1;ram[41][101]=0;ram[41][102]=1;ram[41][103]=1;ram[41][104]=0;ram[41][105]=0;ram[41][106]=1;ram[41][107]=1;ram[41][108]=1;ram[41][109]=1;ram[41][110]=0;ram[41][111]=1;ram[41][112]=1;ram[41][113]=0;ram[41][114]=1;ram[41][115]=1;ram[41][116]=0;ram[41][117]=0;ram[41][118]=1;ram[41][119]=0;ram[41][120]=1;ram[41][121]=0;ram[41][122]=1;ram[41][123]=1;ram[41][124]=0;ram[41][125]=0;ram[41][126]=1;ram[41][127]=1;ram[41][128]=1;ram[41][129]=1;ram[41][130]=0;ram[41][131]=1;ram[41][132]=0;ram[41][133]=0;ram[41][134]=1;ram[41][135]=0;ram[41][136]=0;
        ram[42][0]=1;ram[42][1]=1;ram[42][2]=0;ram[42][3]=0;ram[42][4]=1;ram[42][5]=0;ram[42][6]=1;ram[42][7]=1;ram[42][8]=1;ram[42][9]=1;ram[42][10]=0;ram[42][11]=1;ram[42][12]=1;ram[42][13]=0;ram[42][14]=0;ram[42][15]=1;ram[42][16]=1;ram[42][17]=1;ram[42][18]=1;ram[42][19]=1;ram[42][20]=0;ram[42][21]=0;ram[42][22]=0;ram[42][23]=1;ram[42][24]=0;ram[42][25]=1;ram[42][26]=1;ram[42][27]=0;ram[42][28]=0;ram[42][29]=1;ram[42][30]=1;ram[42][31]=0;ram[42][32]=0;ram[42][33]=1;ram[42][34]=0;ram[42][35]=1;ram[42][36]=0;ram[42][37]=1;ram[42][38]=0;ram[42][39]=1;ram[42][40]=1;ram[42][41]=1;ram[42][42]=0;ram[42][43]=1;ram[42][44]=0;ram[42][45]=0;ram[42][46]=0;ram[42][47]=1;ram[42][48]=1;ram[42][49]=0;ram[42][50]=1;ram[42][51]=1;ram[42][52]=1;ram[42][53]=1;ram[42][54]=1;ram[42][55]=0;ram[42][56]=0;ram[42][57]=1;ram[42][58]=0;ram[42][59]=1;ram[42][60]=1;ram[42][61]=0;ram[42][62]=1;ram[42][63]=0;ram[42][64]=1;ram[42][65]=1;ram[42][66]=1;ram[42][67]=0;ram[42][68]=0;ram[42][69]=1;ram[42][70]=0;ram[42][71]=1;ram[42][72]=1;ram[42][73]=1;ram[42][74]=1;ram[42][75]=1;ram[42][76]=1;ram[42][77]=0;ram[42][78]=1;ram[42][79]=1;ram[42][80]=1;ram[42][81]=1;ram[42][82]=1;ram[42][83]=1;ram[42][84]=1;ram[42][85]=1;ram[42][86]=1;ram[42][87]=1;ram[42][88]=1;ram[42][89]=0;ram[42][90]=1;ram[42][91]=0;ram[42][92]=1;ram[42][93]=1;ram[42][94]=0;ram[42][95]=0;ram[42][96]=0;ram[42][97]=1;ram[42][98]=0;ram[42][99]=1;ram[42][100]=1;ram[42][101]=0;ram[42][102]=0;ram[42][103]=1;ram[42][104]=0;ram[42][105]=1;ram[42][106]=0;ram[42][107]=0;ram[42][108]=0;ram[42][109]=1;ram[42][110]=0;ram[42][111]=0;ram[42][112]=1;ram[42][113]=1;ram[42][114]=1;ram[42][115]=1;ram[42][116]=0;ram[42][117]=1;ram[42][118]=0;ram[42][119]=1;ram[42][120]=0;ram[42][121]=0;ram[42][122]=0;ram[42][123]=1;ram[42][124]=1;ram[42][125]=1;ram[42][126]=1;ram[42][127]=0;ram[42][128]=0;ram[42][129]=0;ram[42][130]=1;ram[42][131]=0;ram[42][132]=0;ram[42][133]=1;ram[42][134]=1;ram[42][135]=0;ram[42][136]=0;
        ram[43][0]=1;ram[43][1]=1;ram[43][2]=1;ram[43][3]=0;ram[43][4]=1;ram[43][5]=1;ram[43][6]=1;ram[43][7]=1;ram[43][8]=0;ram[43][9]=0;ram[43][10]=1;ram[43][11]=0;ram[43][12]=0;ram[43][13]=1;ram[43][14]=0;ram[43][15]=1;ram[43][16]=1;ram[43][17]=0;ram[43][18]=1;ram[43][19]=0;ram[43][20]=1;ram[43][21]=1;ram[43][22]=0;ram[43][23]=1;ram[43][24]=0;ram[43][25]=1;ram[43][26]=1;ram[43][27]=1;ram[43][28]=0;ram[43][29]=1;ram[43][30]=1;ram[43][31]=0;ram[43][32]=1;ram[43][33]=1;ram[43][34]=1;ram[43][35]=0;ram[43][36]=0;ram[43][37]=1;ram[43][38]=0;ram[43][39]=1;ram[43][40]=0;ram[43][41]=0;ram[43][42]=1;ram[43][43]=0;ram[43][44]=0;ram[43][45]=1;ram[43][46]=1;ram[43][47]=1;ram[43][48]=1;ram[43][49]=0;ram[43][50]=0;ram[43][51]=0;ram[43][52]=0;ram[43][53]=1;ram[43][54]=1;ram[43][55]=0;ram[43][56]=1;ram[43][57]=0;ram[43][58]=1;ram[43][59]=0;ram[43][60]=1;ram[43][61]=1;ram[43][62]=1;ram[43][63]=0;ram[43][64]=1;ram[43][65]=1;ram[43][66]=1;ram[43][67]=0;ram[43][68]=1;ram[43][69]=1;ram[43][70]=0;ram[43][71]=1;ram[43][72]=0;ram[43][73]=1;ram[43][74]=1;ram[43][75]=0;ram[43][76]=0;ram[43][77]=1;ram[43][78]=1;ram[43][79]=1;ram[43][80]=1;ram[43][81]=1;ram[43][82]=1;ram[43][83]=1;ram[43][84]=1;ram[43][85]=1;ram[43][86]=1;ram[43][87]=1;ram[43][88]=0;ram[43][89]=0;ram[43][90]=1;ram[43][91]=1;ram[43][92]=1;ram[43][93]=1;ram[43][94]=0;ram[43][95]=0;ram[43][96]=0;ram[43][97]=1;ram[43][98]=1;ram[43][99]=1;ram[43][100]=1;ram[43][101]=1;ram[43][102]=0;ram[43][103]=1;ram[43][104]=0;ram[43][105]=0;ram[43][106]=1;ram[43][107]=0;ram[43][108]=1;ram[43][109]=0;ram[43][110]=1;ram[43][111]=1;ram[43][112]=1;ram[43][113]=0;ram[43][114]=1;ram[43][115]=1;ram[43][116]=1;ram[43][117]=1;ram[43][118]=0;ram[43][119]=1;ram[43][120]=0;ram[43][121]=1;ram[43][122]=0;ram[43][123]=1;ram[43][124]=0;ram[43][125]=1;ram[43][126]=0;ram[43][127]=0;ram[43][128]=1;ram[43][129]=1;ram[43][130]=1;ram[43][131]=0;ram[43][132]=1;ram[43][133]=1;ram[43][134]=0;ram[43][135]=1;ram[43][136]=0;
        ram[44][0]=1;ram[44][1]=1;ram[44][2]=0;ram[44][3]=1;ram[44][4]=1;ram[44][5]=1;ram[44][6]=1;ram[44][7]=0;ram[44][8]=1;ram[44][9]=0;ram[44][10]=1;ram[44][11]=1;ram[44][12]=1;ram[44][13]=0;ram[44][14]=1;ram[44][15]=1;ram[44][16]=1;ram[44][17]=1;ram[44][18]=1;ram[44][19]=1;ram[44][20]=1;ram[44][21]=1;ram[44][22]=0;ram[44][23]=0;ram[44][24]=1;ram[44][25]=1;ram[44][26]=1;ram[44][27]=1;ram[44][28]=1;ram[44][29]=1;ram[44][30]=0;ram[44][31]=1;ram[44][32]=1;ram[44][33]=0;ram[44][34]=0;ram[44][35]=1;ram[44][36]=1;ram[44][37]=1;ram[44][38]=1;ram[44][39]=0;ram[44][40]=1;ram[44][41]=1;ram[44][42]=1;ram[44][43]=0;ram[44][44]=0;ram[44][45]=1;ram[44][46]=1;ram[44][47]=1;ram[44][48]=1;ram[44][49]=1;ram[44][50]=1;ram[44][51]=1;ram[44][52]=1;ram[44][53]=0;ram[44][54]=1;ram[44][55]=1;ram[44][56]=0;ram[44][57]=0;ram[44][58]=1;ram[44][59]=1;ram[44][60]=0;ram[44][61]=0;ram[44][62]=1;ram[44][63]=1;ram[44][64]=1;ram[44][65]=1;ram[44][66]=1;ram[44][67]=0;ram[44][68]=1;ram[44][69]=1;ram[44][70]=1;ram[44][71]=1;ram[44][72]=0;ram[44][73]=1;ram[44][74]=0;ram[44][75]=1;ram[44][76]=0;ram[44][77]=1;ram[44][78]=0;ram[44][79]=1;ram[44][80]=0;ram[44][81]=1;ram[44][82]=0;ram[44][83]=1;ram[44][84]=1;ram[44][85]=0;ram[44][86]=0;ram[44][87]=0;ram[44][88]=0;ram[44][89]=0;ram[44][90]=0;ram[44][91]=1;ram[44][92]=1;ram[44][93]=1;ram[44][94]=0;ram[44][95]=0;ram[44][96]=1;ram[44][97]=0;ram[44][98]=1;ram[44][99]=0;ram[44][100]=0;ram[44][101]=1;ram[44][102]=0;ram[44][103]=1;ram[44][104]=1;ram[44][105]=1;ram[44][106]=0;ram[44][107]=0;ram[44][108]=0;ram[44][109]=1;ram[44][110]=1;ram[44][111]=1;ram[44][112]=1;ram[44][113]=1;ram[44][114]=1;ram[44][115]=0;ram[44][116]=0;ram[44][117]=0;ram[44][118]=1;ram[44][119]=1;ram[44][120]=1;ram[44][121]=1;ram[44][122]=1;ram[44][123]=1;ram[44][124]=1;ram[44][125]=1;ram[44][126]=1;ram[44][127]=0;ram[44][128]=1;ram[44][129]=0;ram[44][130]=1;ram[44][131]=0;ram[44][132]=1;ram[44][133]=1;ram[44][134]=1;ram[44][135]=1;ram[44][136]=0;
        ram[45][0]=0;ram[45][1]=1;ram[45][2]=1;ram[45][3]=0;ram[45][4]=1;ram[45][5]=1;ram[45][6]=1;ram[45][7]=1;ram[45][8]=1;ram[45][9]=1;ram[45][10]=0;ram[45][11]=1;ram[45][12]=1;ram[45][13]=1;ram[45][14]=1;ram[45][15]=1;ram[45][16]=1;ram[45][17]=0;ram[45][18]=1;ram[45][19]=1;ram[45][20]=1;ram[45][21]=1;ram[45][22]=1;ram[45][23]=0;ram[45][24]=1;ram[45][25]=1;ram[45][26]=1;ram[45][27]=1;ram[45][28]=0;ram[45][29]=1;ram[45][30]=1;ram[45][31]=1;ram[45][32]=0;ram[45][33]=1;ram[45][34]=1;ram[45][35]=0;ram[45][36]=1;ram[45][37]=1;ram[45][38]=0;ram[45][39]=0;ram[45][40]=1;ram[45][41]=1;ram[45][42]=1;ram[45][43]=1;ram[45][44]=0;ram[45][45]=0;ram[45][46]=1;ram[45][47]=0;ram[45][48]=1;ram[45][49]=1;ram[45][50]=1;ram[45][51]=1;ram[45][52]=1;ram[45][53]=0;ram[45][54]=1;ram[45][55]=0;ram[45][56]=1;ram[45][57]=1;ram[45][58]=1;ram[45][59]=1;ram[45][60]=0;ram[45][61]=1;ram[45][62]=1;ram[45][63]=1;ram[45][64]=1;ram[45][65]=1;ram[45][66]=1;ram[45][67]=0;ram[45][68]=1;ram[45][69]=0;ram[45][70]=1;ram[45][71]=1;ram[45][72]=1;ram[45][73]=0;ram[45][74]=0;ram[45][75]=1;ram[45][76]=0;ram[45][77]=1;ram[45][78]=0;ram[45][79]=0;ram[45][80]=1;ram[45][81]=0;ram[45][82]=1;ram[45][83]=0;ram[45][84]=1;ram[45][85]=0;ram[45][86]=0;ram[45][87]=1;ram[45][88]=0;ram[45][89]=1;ram[45][90]=0;ram[45][91]=0;ram[45][92]=1;ram[45][93]=0;ram[45][94]=0;ram[45][95]=1;ram[45][96]=1;ram[45][97]=0;ram[45][98]=0;ram[45][99]=0;ram[45][100]=1;ram[45][101]=0;ram[45][102]=1;ram[45][103]=0;ram[45][104]=0;ram[45][105]=0;ram[45][106]=1;ram[45][107]=0;ram[45][108]=0;ram[45][109]=0;ram[45][110]=1;ram[45][111]=1;ram[45][112]=0;ram[45][113]=1;ram[45][114]=0;ram[45][115]=0;ram[45][116]=0;ram[45][117]=1;ram[45][118]=1;ram[45][119]=0;ram[45][120]=1;ram[45][121]=0;ram[45][122]=1;ram[45][123]=1;ram[45][124]=1;ram[45][125]=0;ram[45][126]=0;ram[45][127]=1;ram[45][128]=0;ram[45][129]=1;ram[45][130]=1;ram[45][131]=1;ram[45][132]=1;ram[45][133]=1;ram[45][134]=0;ram[45][135]=0;ram[45][136]=0;
        ram[46][0]=1;ram[46][1]=0;ram[46][2]=1;ram[46][3]=1;ram[46][4]=0;ram[46][5]=1;ram[46][6]=1;ram[46][7]=0;ram[46][8]=0;ram[46][9]=0;ram[46][10]=1;ram[46][11]=1;ram[46][12]=1;ram[46][13]=0;ram[46][14]=1;ram[46][15]=0;ram[46][16]=1;ram[46][17]=1;ram[46][18]=1;ram[46][19]=0;ram[46][20]=0;ram[46][21]=0;ram[46][22]=0;ram[46][23]=1;ram[46][24]=1;ram[46][25]=0;ram[46][26]=1;ram[46][27]=1;ram[46][28]=0;ram[46][29]=1;ram[46][30]=0;ram[46][31]=1;ram[46][32]=1;ram[46][33]=1;ram[46][34]=1;ram[46][35]=0;ram[46][36]=1;ram[46][37]=1;ram[46][38]=0;ram[46][39]=0;ram[46][40]=1;ram[46][41]=1;ram[46][42]=0;ram[46][43]=1;ram[46][44]=1;ram[46][45]=1;ram[46][46]=1;ram[46][47]=1;ram[46][48]=0;ram[46][49]=1;ram[46][50]=1;ram[46][51]=0;ram[46][52]=0;ram[46][53]=1;ram[46][54]=1;ram[46][55]=0;ram[46][56]=1;ram[46][57]=1;ram[46][58]=1;ram[46][59]=1;ram[46][60]=1;ram[46][61]=1;ram[46][62]=1;ram[46][63]=1;ram[46][64]=1;ram[46][65]=0;ram[46][66]=0;ram[46][67]=1;ram[46][68]=1;ram[46][69]=0;ram[46][70]=1;ram[46][71]=1;ram[46][72]=0;ram[46][73]=0;ram[46][74]=0;ram[46][75]=1;ram[46][76]=0;ram[46][77]=1;ram[46][78]=1;ram[46][79]=1;ram[46][80]=0;ram[46][81]=1;ram[46][82]=0;ram[46][83]=1;ram[46][84]=0;ram[46][85]=1;ram[46][86]=1;ram[46][87]=1;ram[46][88]=0;ram[46][89]=1;ram[46][90]=1;ram[46][91]=0;ram[46][92]=0;ram[46][93]=0;ram[46][94]=1;ram[46][95]=0;ram[46][96]=1;ram[46][97]=0;ram[46][98]=1;ram[46][99]=0;ram[46][100]=0;ram[46][101]=1;ram[46][102]=1;ram[46][103]=1;ram[46][104]=1;ram[46][105]=1;ram[46][106]=0;ram[46][107]=0;ram[46][108]=0;ram[46][109]=0;ram[46][110]=0;ram[46][111]=0;ram[46][112]=0;ram[46][113]=0;ram[46][114]=0;ram[46][115]=1;ram[46][116]=1;ram[46][117]=1;ram[46][118]=1;ram[46][119]=0;ram[46][120]=1;ram[46][121]=0;ram[46][122]=1;ram[46][123]=1;ram[46][124]=0;ram[46][125]=1;ram[46][126]=0;ram[46][127]=0;ram[46][128]=0;ram[46][129]=1;ram[46][130]=1;ram[46][131]=1;ram[46][132]=0;ram[46][133]=1;ram[46][134]=0;ram[46][135]=1;ram[46][136]=1;
        ram[47][0]=0;ram[47][1]=1;ram[47][2]=0;ram[47][3]=1;ram[47][4]=0;ram[47][5]=0;ram[47][6]=1;ram[47][7]=1;ram[47][8]=1;ram[47][9]=1;ram[47][10]=0;ram[47][11]=1;ram[47][12]=0;ram[47][13]=1;ram[47][14]=1;ram[47][15]=1;ram[47][16]=0;ram[47][17]=1;ram[47][18]=1;ram[47][19]=1;ram[47][20]=1;ram[47][21]=0;ram[47][22]=0;ram[47][23]=1;ram[47][24]=0;ram[47][25]=0;ram[47][26]=1;ram[47][27]=0;ram[47][28]=1;ram[47][29]=0;ram[47][30]=1;ram[47][31]=1;ram[47][32]=0;ram[47][33]=1;ram[47][34]=0;ram[47][35]=1;ram[47][36]=1;ram[47][37]=0;ram[47][38]=0;ram[47][39]=1;ram[47][40]=0;ram[47][41]=1;ram[47][42]=1;ram[47][43]=1;ram[47][44]=1;ram[47][45]=0;ram[47][46]=1;ram[47][47]=1;ram[47][48]=1;ram[47][49]=0;ram[47][50]=1;ram[47][51]=0;ram[47][52]=1;ram[47][53]=0;ram[47][54]=1;ram[47][55]=1;ram[47][56]=1;ram[47][57]=1;ram[47][58]=0;ram[47][59]=1;ram[47][60]=0;ram[47][61]=0;ram[47][62]=0;ram[47][63]=1;ram[47][64]=1;ram[47][65]=1;ram[47][66]=1;ram[47][67]=1;ram[47][68]=1;ram[47][69]=1;ram[47][70]=1;ram[47][71]=1;ram[47][72]=1;ram[47][73]=1;ram[47][74]=1;ram[47][75]=1;ram[47][76]=1;ram[47][77]=0;ram[47][78]=1;ram[47][79]=1;ram[47][80]=0;ram[47][81]=1;ram[47][82]=0;ram[47][83]=0;ram[47][84]=1;ram[47][85]=1;ram[47][86]=1;ram[47][87]=1;ram[47][88]=0;ram[47][89]=1;ram[47][90]=1;ram[47][91]=0;ram[47][92]=1;ram[47][93]=0;ram[47][94]=1;ram[47][95]=1;ram[47][96]=0;ram[47][97]=1;ram[47][98]=0;ram[47][99]=0;ram[47][100]=1;ram[47][101]=1;ram[47][102]=0;ram[47][103]=1;ram[47][104]=1;ram[47][105]=1;ram[47][106]=0;ram[47][107]=1;ram[47][108]=1;ram[47][109]=1;ram[47][110]=1;ram[47][111]=1;ram[47][112]=0;ram[47][113]=0;ram[47][114]=1;ram[47][115]=1;ram[47][116]=1;ram[47][117]=0;ram[47][118]=1;ram[47][119]=1;ram[47][120]=1;ram[47][121]=1;ram[47][122]=1;ram[47][123]=1;ram[47][124]=0;ram[47][125]=1;ram[47][126]=1;ram[47][127]=1;ram[47][128]=0;ram[47][129]=1;ram[47][130]=1;ram[47][131]=1;ram[47][132]=1;ram[47][133]=0;ram[47][134]=1;ram[47][135]=1;ram[47][136]=0;
        ram[48][0]=1;ram[48][1]=1;ram[48][2]=1;ram[48][3]=0;ram[48][4]=1;ram[48][5]=0;ram[48][6]=1;ram[48][7]=0;ram[48][8]=1;ram[48][9]=0;ram[48][10]=1;ram[48][11]=1;ram[48][12]=0;ram[48][13]=0;ram[48][14]=1;ram[48][15]=0;ram[48][16]=1;ram[48][17]=1;ram[48][18]=1;ram[48][19]=1;ram[48][20]=1;ram[48][21]=0;ram[48][22]=1;ram[48][23]=0;ram[48][24]=1;ram[48][25]=1;ram[48][26]=1;ram[48][27]=1;ram[48][28]=1;ram[48][29]=1;ram[48][30]=1;ram[48][31]=1;ram[48][32]=1;ram[48][33]=1;ram[48][34]=1;ram[48][35]=1;ram[48][36]=1;ram[48][37]=0;ram[48][38]=0;ram[48][39]=0;ram[48][40]=0;ram[48][41]=1;ram[48][42]=1;ram[48][43]=1;ram[48][44]=1;ram[48][45]=0;ram[48][46]=1;ram[48][47]=0;ram[48][48]=1;ram[48][49]=0;ram[48][50]=1;ram[48][51]=1;ram[48][52]=1;ram[48][53]=1;ram[48][54]=0;ram[48][55]=1;ram[48][56]=0;ram[48][57]=1;ram[48][58]=0;ram[48][59]=0;ram[48][60]=0;ram[48][61]=1;ram[48][62]=1;ram[48][63]=1;ram[48][64]=1;ram[48][65]=0;ram[48][66]=0;ram[48][67]=1;ram[48][68]=1;ram[48][69]=0;ram[48][70]=0;ram[48][71]=1;ram[48][72]=1;ram[48][73]=1;ram[48][74]=1;ram[48][75]=1;ram[48][76]=0;ram[48][77]=1;ram[48][78]=1;ram[48][79]=1;ram[48][80]=1;ram[48][81]=1;ram[48][82]=1;ram[48][83]=0;ram[48][84]=1;ram[48][85]=1;ram[48][86]=0;ram[48][87]=1;ram[48][88]=1;ram[48][89]=1;ram[48][90]=0;ram[48][91]=0;ram[48][92]=1;ram[48][93]=0;ram[48][94]=1;ram[48][95]=1;ram[48][96]=1;ram[48][97]=1;ram[48][98]=1;ram[48][99]=0;ram[48][100]=1;ram[48][101]=0;ram[48][102]=1;ram[48][103]=1;ram[48][104]=1;ram[48][105]=1;ram[48][106]=1;ram[48][107]=0;ram[48][108]=1;ram[48][109]=0;ram[48][110]=0;ram[48][111]=1;ram[48][112]=1;ram[48][113]=1;ram[48][114]=1;ram[48][115]=1;ram[48][116]=1;ram[48][117]=1;ram[48][118]=1;ram[48][119]=0;ram[48][120]=1;ram[48][121]=0;ram[48][122]=1;ram[48][123]=0;ram[48][124]=0;ram[48][125]=0;ram[48][126]=1;ram[48][127]=1;ram[48][128]=1;ram[48][129]=1;ram[48][130]=0;ram[48][131]=1;ram[48][132]=1;ram[48][133]=1;ram[48][134]=0;ram[48][135]=0;ram[48][136]=0;
        ram[49][0]=0;ram[49][1]=0;ram[49][2]=1;ram[49][3]=1;ram[49][4]=1;ram[49][5]=1;ram[49][6]=1;ram[49][7]=1;ram[49][8]=1;ram[49][9]=1;ram[49][10]=1;ram[49][11]=0;ram[49][12]=0;ram[49][13]=1;ram[49][14]=0;ram[49][15]=0;ram[49][16]=1;ram[49][17]=0;ram[49][18]=1;ram[49][19]=1;ram[49][20]=1;ram[49][21]=1;ram[49][22]=0;ram[49][23]=1;ram[49][24]=1;ram[49][25]=1;ram[49][26]=0;ram[49][27]=1;ram[49][28]=0;ram[49][29]=1;ram[49][30]=1;ram[49][31]=1;ram[49][32]=0;ram[49][33]=0;ram[49][34]=0;ram[49][35]=1;ram[49][36]=1;ram[49][37]=0;ram[49][38]=1;ram[49][39]=0;ram[49][40]=1;ram[49][41]=1;ram[49][42]=0;ram[49][43]=1;ram[49][44]=1;ram[49][45]=1;ram[49][46]=0;ram[49][47]=1;ram[49][48]=1;ram[49][49]=0;ram[49][50]=1;ram[49][51]=0;ram[49][52]=1;ram[49][53]=1;ram[49][54]=1;ram[49][55]=0;ram[49][56]=1;ram[49][57]=0;ram[49][58]=1;ram[49][59]=0;ram[49][60]=0;ram[49][61]=1;ram[49][62]=0;ram[49][63]=1;ram[49][64]=1;ram[49][65]=1;ram[49][66]=0;ram[49][67]=0;ram[49][68]=1;ram[49][69]=1;ram[49][70]=1;ram[49][71]=0;ram[49][72]=1;ram[49][73]=1;ram[49][74]=0;ram[49][75]=1;ram[49][76]=0;ram[49][77]=1;ram[49][78]=1;ram[49][79]=0;ram[49][80]=1;ram[49][81]=1;ram[49][82]=1;ram[49][83]=1;ram[49][84]=1;ram[49][85]=1;ram[49][86]=0;ram[49][87]=0;ram[49][88]=0;ram[49][89]=1;ram[49][90]=0;ram[49][91]=0;ram[49][92]=0;ram[49][93]=1;ram[49][94]=1;ram[49][95]=0;ram[49][96]=0;ram[49][97]=0;ram[49][98]=0;ram[49][99]=0;ram[49][100]=0;ram[49][101]=1;ram[49][102]=1;ram[49][103]=1;ram[49][104]=0;ram[49][105]=1;ram[49][106]=0;ram[49][107]=1;ram[49][108]=1;ram[49][109]=1;ram[49][110]=1;ram[49][111]=0;ram[49][112]=1;ram[49][113]=1;ram[49][114]=1;ram[49][115]=0;ram[49][116]=0;ram[49][117]=1;ram[49][118]=0;ram[49][119]=0;ram[49][120]=1;ram[49][121]=0;ram[49][122]=0;ram[49][123]=0;ram[49][124]=1;ram[49][125]=1;ram[49][126]=1;ram[49][127]=1;ram[49][128]=1;ram[49][129]=0;ram[49][130]=1;ram[49][131]=1;ram[49][132]=1;ram[49][133]=1;ram[49][134]=0;ram[49][135]=1;ram[49][136]=1;
        ram[50][0]=1;ram[50][1]=0;ram[50][2]=1;ram[50][3]=1;ram[50][4]=1;ram[50][5]=1;ram[50][6]=0;ram[50][7]=0;ram[50][8]=1;ram[50][9]=1;ram[50][10]=1;ram[50][11]=1;ram[50][12]=0;ram[50][13]=0;ram[50][14]=0;ram[50][15]=1;ram[50][16]=1;ram[50][17]=0;ram[50][18]=0;ram[50][19]=1;ram[50][20]=0;ram[50][21]=0;ram[50][22]=1;ram[50][23]=1;ram[50][24]=1;ram[50][25]=1;ram[50][26]=1;ram[50][27]=1;ram[50][28]=0;ram[50][29]=1;ram[50][30]=1;ram[50][31]=1;ram[50][32]=1;ram[50][33]=1;ram[50][34]=0;ram[50][35]=0;ram[50][36]=1;ram[50][37]=1;ram[50][38]=0;ram[50][39]=1;ram[50][40]=0;ram[50][41]=1;ram[50][42]=0;ram[50][43]=0;ram[50][44]=0;ram[50][45]=1;ram[50][46]=0;ram[50][47]=1;ram[50][48]=1;ram[50][49]=0;ram[50][50]=1;ram[50][51]=1;ram[50][52]=0;ram[50][53]=1;ram[50][54]=1;ram[50][55]=1;ram[50][56]=1;ram[50][57]=0;ram[50][58]=1;ram[50][59]=0;ram[50][60]=1;ram[50][61]=1;ram[50][62]=1;ram[50][63]=1;ram[50][64]=0;ram[50][65]=1;ram[50][66]=0;ram[50][67]=0;ram[50][68]=1;ram[50][69]=0;ram[50][70]=1;ram[50][71]=1;ram[50][72]=0;ram[50][73]=0;ram[50][74]=0;ram[50][75]=1;ram[50][76]=0;ram[50][77]=1;ram[50][78]=0;ram[50][79]=0;ram[50][80]=0;ram[50][81]=0;ram[50][82]=0;ram[50][83]=0;ram[50][84]=1;ram[50][85]=1;ram[50][86]=0;ram[50][87]=0;ram[50][88]=1;ram[50][89]=1;ram[50][90]=0;ram[50][91]=1;ram[50][92]=0;ram[50][93]=1;ram[50][94]=1;ram[50][95]=1;ram[50][96]=0;ram[50][97]=1;ram[50][98]=1;ram[50][99]=0;ram[50][100]=1;ram[50][101]=1;ram[50][102]=0;ram[50][103]=1;ram[50][104]=1;ram[50][105]=1;ram[50][106]=0;ram[50][107]=1;ram[50][108]=1;ram[50][109]=1;ram[50][110]=1;ram[50][111]=1;ram[50][112]=1;ram[50][113]=1;ram[50][114]=1;ram[50][115]=1;ram[50][116]=0;ram[50][117]=1;ram[50][118]=1;ram[50][119]=1;ram[50][120]=1;ram[50][121]=0;ram[50][122]=0;ram[50][123]=1;ram[50][124]=0;ram[50][125]=1;ram[50][126]=1;ram[50][127]=1;ram[50][128]=1;ram[50][129]=1;ram[50][130]=0;ram[50][131]=1;ram[50][132]=1;ram[50][133]=1;ram[50][134]=0;ram[50][135]=1;ram[50][136]=1;
        ram[51][0]=1;ram[51][1]=1;ram[51][2]=1;ram[51][3]=0;ram[51][4]=1;ram[51][5]=1;ram[51][6]=0;ram[51][7]=1;ram[51][8]=0;ram[51][9]=0;ram[51][10]=1;ram[51][11]=0;ram[51][12]=0;ram[51][13]=1;ram[51][14]=0;ram[51][15]=0;ram[51][16]=1;ram[51][17]=1;ram[51][18]=1;ram[51][19]=0;ram[51][20]=1;ram[51][21]=1;ram[51][22]=1;ram[51][23]=1;ram[51][24]=1;ram[51][25]=0;ram[51][26]=1;ram[51][27]=1;ram[51][28]=1;ram[51][29]=0;ram[51][30]=0;ram[51][31]=0;ram[51][32]=0;ram[51][33]=0;ram[51][34]=0;ram[51][35]=0;ram[51][36]=1;ram[51][37]=0;ram[51][38]=0;ram[51][39]=1;ram[51][40]=1;ram[51][41]=1;ram[51][42]=1;ram[51][43]=1;ram[51][44]=1;ram[51][45]=1;ram[51][46]=1;ram[51][47]=0;ram[51][48]=0;ram[51][49]=0;ram[51][50]=1;ram[51][51]=0;ram[51][52]=0;ram[51][53]=1;ram[51][54]=1;ram[51][55]=1;ram[51][56]=1;ram[51][57]=1;ram[51][58]=0;ram[51][59]=0;ram[51][60]=1;ram[51][61]=1;ram[51][62]=1;ram[51][63]=1;ram[51][64]=0;ram[51][65]=1;ram[51][66]=0;ram[51][67]=1;ram[51][68]=1;ram[51][69]=0;ram[51][70]=1;ram[51][71]=1;ram[51][72]=0;ram[51][73]=1;ram[51][74]=0;ram[51][75]=1;ram[51][76]=0;ram[51][77]=1;ram[51][78]=1;ram[51][79]=1;ram[51][80]=0;ram[51][81]=1;ram[51][82]=0;ram[51][83]=0;ram[51][84]=1;ram[51][85]=1;ram[51][86]=0;ram[51][87]=0;ram[51][88]=1;ram[51][89]=1;ram[51][90]=1;ram[51][91]=1;ram[51][92]=1;ram[51][93]=0;ram[51][94]=0;ram[51][95]=1;ram[51][96]=1;ram[51][97]=1;ram[51][98]=1;ram[51][99]=1;ram[51][100]=1;ram[51][101]=0;ram[51][102]=1;ram[51][103]=0;ram[51][104]=0;ram[51][105]=0;ram[51][106]=1;ram[51][107]=0;ram[51][108]=1;ram[51][109]=1;ram[51][110]=1;ram[51][111]=0;ram[51][112]=1;ram[51][113]=1;ram[51][114]=1;ram[51][115]=1;ram[51][116]=0;ram[51][117]=1;ram[51][118]=1;ram[51][119]=0;ram[51][120]=1;ram[51][121]=1;ram[51][122]=0;ram[51][123]=1;ram[51][124]=1;ram[51][125]=1;ram[51][126]=0;ram[51][127]=0;ram[51][128]=1;ram[51][129]=1;ram[51][130]=1;ram[51][131]=0;ram[51][132]=0;ram[51][133]=1;ram[51][134]=1;ram[51][135]=1;ram[51][136]=1;
        ram[52][0]=1;ram[52][1]=0;ram[52][2]=1;ram[52][3]=0;ram[52][4]=0;ram[52][5]=1;ram[52][6]=0;ram[52][7]=0;ram[52][8]=0;ram[52][9]=1;ram[52][10]=1;ram[52][11]=1;ram[52][12]=1;ram[52][13]=0;ram[52][14]=1;ram[52][15]=1;ram[52][16]=0;ram[52][17]=0;ram[52][18]=1;ram[52][19]=0;ram[52][20]=0;ram[52][21]=1;ram[52][22]=1;ram[52][23]=1;ram[52][24]=0;ram[52][25]=0;ram[52][26]=1;ram[52][27]=0;ram[52][28]=1;ram[52][29]=0;ram[52][30]=0;ram[52][31]=1;ram[52][32]=1;ram[52][33]=1;ram[52][34]=0;ram[52][35]=1;ram[52][36]=0;ram[52][37]=0;ram[52][38]=0;ram[52][39]=1;ram[52][40]=1;ram[52][41]=1;ram[52][42]=1;ram[52][43]=1;ram[52][44]=1;ram[52][45]=1;ram[52][46]=0;ram[52][47]=0;ram[52][48]=1;ram[52][49]=0;ram[52][50]=1;ram[52][51]=0;ram[52][52]=0;ram[52][53]=0;ram[52][54]=0;ram[52][55]=1;ram[52][56]=1;ram[52][57]=1;ram[52][58]=1;ram[52][59]=1;ram[52][60]=1;ram[52][61]=1;ram[52][62]=1;ram[52][63]=0;ram[52][64]=1;ram[52][65]=1;ram[52][66]=0;ram[52][67]=0;ram[52][68]=1;ram[52][69]=0;ram[52][70]=0;ram[52][71]=0;ram[52][72]=1;ram[52][73]=0;ram[52][74]=1;ram[52][75]=0;ram[52][76]=1;ram[52][77]=0;ram[52][78]=0;ram[52][79]=0;ram[52][80]=0;ram[52][81]=0;ram[52][82]=1;ram[52][83]=1;ram[52][84]=1;ram[52][85]=1;ram[52][86]=0;ram[52][87]=1;ram[52][88]=0;ram[52][89]=0;ram[52][90]=1;ram[52][91]=1;ram[52][92]=0;ram[52][93]=1;ram[52][94]=1;ram[52][95]=1;ram[52][96]=1;ram[52][97]=0;ram[52][98]=0;ram[52][99]=1;ram[52][100]=0;ram[52][101]=0;ram[52][102]=1;ram[52][103]=1;ram[52][104]=0;ram[52][105]=1;ram[52][106]=1;ram[52][107]=0;ram[52][108]=1;ram[52][109]=1;ram[52][110]=0;ram[52][111]=1;ram[52][112]=0;ram[52][113]=0;ram[52][114]=1;ram[52][115]=1;ram[52][116]=0;ram[52][117]=1;ram[52][118]=0;ram[52][119]=1;ram[52][120]=1;ram[52][121]=1;ram[52][122]=1;ram[52][123]=1;ram[52][124]=1;ram[52][125]=1;ram[52][126]=0;ram[52][127]=1;ram[52][128]=1;ram[52][129]=1;ram[52][130]=1;ram[52][131]=1;ram[52][132]=1;ram[52][133]=1;ram[52][134]=1;ram[52][135]=1;ram[52][136]=1;
        ram[53][0]=1;ram[53][1]=1;ram[53][2]=0;ram[53][3]=1;ram[53][4]=1;ram[53][5]=0;ram[53][6]=1;ram[53][7]=0;ram[53][8]=1;ram[53][9]=1;ram[53][10]=1;ram[53][11]=1;ram[53][12]=1;ram[53][13]=1;ram[53][14]=1;ram[53][15]=1;ram[53][16]=1;ram[53][17]=1;ram[53][18]=1;ram[53][19]=1;ram[53][20]=1;ram[53][21]=1;ram[53][22]=1;ram[53][23]=0;ram[53][24]=1;ram[53][25]=0;ram[53][26]=1;ram[53][27]=0;ram[53][28]=1;ram[53][29]=1;ram[53][30]=1;ram[53][31]=1;ram[53][32]=1;ram[53][33]=1;ram[53][34]=1;ram[53][35]=0;ram[53][36]=0;ram[53][37]=0;ram[53][38]=0;ram[53][39]=1;ram[53][40]=1;ram[53][41]=1;ram[53][42]=0;ram[53][43]=1;ram[53][44]=1;ram[53][45]=0;ram[53][46]=1;ram[53][47]=0;ram[53][48]=1;ram[53][49]=1;ram[53][50]=1;ram[53][51]=0;ram[53][52]=0;ram[53][53]=1;ram[53][54]=1;ram[53][55]=1;ram[53][56]=0;ram[53][57]=0;ram[53][58]=1;ram[53][59]=1;ram[53][60]=1;ram[53][61]=1;ram[53][62]=0;ram[53][63]=1;ram[53][64]=1;ram[53][65]=1;ram[53][66]=0;ram[53][67]=1;ram[53][68]=0;ram[53][69]=1;ram[53][70]=1;ram[53][71]=0;ram[53][72]=0;ram[53][73]=0;ram[53][74]=1;ram[53][75]=1;ram[53][76]=1;ram[53][77]=1;ram[53][78]=1;ram[53][79]=1;ram[53][80]=1;ram[53][81]=1;ram[53][82]=1;ram[53][83]=0;ram[53][84]=0;ram[53][85]=1;ram[53][86]=1;ram[53][87]=0;ram[53][88]=1;ram[53][89]=0;ram[53][90]=1;ram[53][91]=1;ram[53][92]=1;ram[53][93]=0;ram[53][94]=0;ram[53][95]=0;ram[53][96]=0;ram[53][97]=1;ram[53][98]=1;ram[53][99]=0;ram[53][100]=1;ram[53][101]=1;ram[53][102]=1;ram[53][103]=1;ram[53][104]=1;ram[53][105]=0;ram[53][106]=1;ram[53][107]=1;ram[53][108]=1;ram[53][109]=1;ram[53][110]=0;ram[53][111]=1;ram[53][112]=1;ram[53][113]=1;ram[53][114]=1;ram[53][115]=1;ram[53][116]=1;ram[53][117]=1;ram[53][118]=1;ram[53][119]=1;ram[53][120]=1;ram[53][121]=1;ram[53][122]=1;ram[53][123]=0;ram[53][124]=1;ram[53][125]=1;ram[53][126]=1;ram[53][127]=1;ram[53][128]=0;ram[53][129]=1;ram[53][130]=0;ram[53][131]=1;ram[53][132]=1;ram[53][133]=0;ram[53][134]=0;ram[53][135]=1;ram[53][136]=1;
        ram[54][0]=0;ram[54][1]=1;ram[54][2]=1;ram[54][3]=0;ram[54][4]=1;ram[54][5]=0;ram[54][6]=0;ram[54][7]=1;ram[54][8]=1;ram[54][9]=1;ram[54][10]=0;ram[54][11]=1;ram[54][12]=0;ram[54][13]=0;ram[54][14]=1;ram[54][15]=0;ram[54][16]=1;ram[54][17]=0;ram[54][18]=1;ram[54][19]=1;ram[54][20]=0;ram[54][21]=1;ram[54][22]=0;ram[54][23]=1;ram[54][24]=1;ram[54][25]=1;ram[54][26]=1;ram[54][27]=0;ram[54][28]=1;ram[54][29]=1;ram[54][30]=0;ram[54][31]=1;ram[54][32]=0;ram[54][33]=1;ram[54][34]=1;ram[54][35]=1;ram[54][36]=0;ram[54][37]=0;ram[54][38]=1;ram[54][39]=1;ram[54][40]=1;ram[54][41]=1;ram[54][42]=1;ram[54][43]=1;ram[54][44]=1;ram[54][45]=1;ram[54][46]=0;ram[54][47]=1;ram[54][48]=1;ram[54][49]=0;ram[54][50]=1;ram[54][51]=0;ram[54][52]=0;ram[54][53]=1;ram[54][54]=1;ram[54][55]=1;ram[54][56]=1;ram[54][57]=1;ram[54][58]=1;ram[54][59]=0;ram[54][60]=1;ram[54][61]=1;ram[54][62]=0;ram[54][63]=1;ram[54][64]=1;ram[54][65]=1;ram[54][66]=1;ram[54][67]=0;ram[54][68]=1;ram[54][69]=1;ram[54][70]=0;ram[54][71]=0;ram[54][72]=1;ram[54][73]=1;ram[54][74]=1;ram[54][75]=0;ram[54][76]=1;ram[54][77]=1;ram[54][78]=1;ram[54][79]=1;ram[54][80]=1;ram[54][81]=1;ram[54][82]=1;ram[54][83]=1;ram[54][84]=0;ram[54][85]=1;ram[54][86]=1;ram[54][87]=1;ram[54][88]=0;ram[54][89]=1;ram[54][90]=1;ram[54][91]=1;ram[54][92]=1;ram[54][93]=0;ram[54][94]=1;ram[54][95]=0;ram[54][96]=0;ram[54][97]=1;ram[54][98]=1;ram[54][99]=0;ram[54][100]=1;ram[54][101]=0;ram[54][102]=1;ram[54][103]=0;ram[54][104]=1;ram[54][105]=1;ram[54][106]=0;ram[54][107]=0;ram[54][108]=1;ram[54][109]=1;ram[54][110]=1;ram[54][111]=0;ram[54][112]=1;ram[54][113]=0;ram[54][114]=0;ram[54][115]=1;ram[54][116]=1;ram[54][117]=1;ram[54][118]=1;ram[54][119]=0;ram[54][120]=1;ram[54][121]=0;ram[54][122]=1;ram[54][123]=1;ram[54][124]=0;ram[54][125]=1;ram[54][126]=1;ram[54][127]=1;ram[54][128]=0;ram[54][129]=1;ram[54][130]=0;ram[54][131]=0;ram[54][132]=0;ram[54][133]=0;ram[54][134]=1;ram[54][135]=0;ram[54][136]=0;
        ram[55][0]=0;ram[55][1]=0;ram[55][2]=0;ram[55][3]=1;ram[55][4]=1;ram[55][5]=1;ram[55][6]=1;ram[55][7]=1;ram[55][8]=0;ram[55][9]=1;ram[55][10]=1;ram[55][11]=1;ram[55][12]=1;ram[55][13]=1;ram[55][14]=1;ram[55][15]=0;ram[55][16]=1;ram[55][17]=1;ram[55][18]=1;ram[55][19]=1;ram[55][20]=1;ram[55][21]=0;ram[55][22]=0;ram[55][23]=1;ram[55][24]=0;ram[55][25]=1;ram[55][26]=1;ram[55][27]=1;ram[55][28]=1;ram[55][29]=1;ram[55][30]=0;ram[55][31]=1;ram[55][32]=1;ram[55][33]=1;ram[55][34]=0;ram[55][35]=1;ram[55][36]=1;ram[55][37]=1;ram[55][38]=0;ram[55][39]=1;ram[55][40]=1;ram[55][41]=1;ram[55][42]=1;ram[55][43]=1;ram[55][44]=1;ram[55][45]=0;ram[55][46]=1;ram[55][47]=1;ram[55][48]=1;ram[55][49]=1;ram[55][50]=1;ram[55][51]=0;ram[55][52]=1;ram[55][53]=1;ram[55][54]=1;ram[55][55]=1;ram[55][56]=1;ram[55][57]=0;ram[55][58]=1;ram[55][59]=0;ram[55][60]=1;ram[55][61]=0;ram[55][62]=1;ram[55][63]=1;ram[55][64]=0;ram[55][65]=1;ram[55][66]=0;ram[55][67]=0;ram[55][68]=1;ram[55][69]=1;ram[55][70]=1;ram[55][71]=1;ram[55][72]=0;ram[55][73]=0;ram[55][74]=0;ram[55][75]=0;ram[55][76]=1;ram[55][77]=1;ram[55][78]=1;ram[55][79]=1;ram[55][80]=1;ram[55][81]=0;ram[55][82]=0;ram[55][83]=0;ram[55][84]=1;ram[55][85]=1;ram[55][86]=0;ram[55][87]=1;ram[55][88]=0;ram[55][89]=1;ram[55][90]=0;ram[55][91]=0;ram[55][92]=1;ram[55][93]=1;ram[55][94]=1;ram[55][95]=1;ram[55][96]=1;ram[55][97]=1;ram[55][98]=1;ram[55][99]=1;ram[55][100]=1;ram[55][101]=1;ram[55][102]=1;ram[55][103]=1;ram[55][104]=0;ram[55][105]=0;ram[55][106]=0;ram[55][107]=0;ram[55][108]=1;ram[55][109]=0;ram[55][110]=1;ram[55][111]=1;ram[55][112]=1;ram[55][113]=1;ram[55][114]=1;ram[55][115]=1;ram[55][116]=1;ram[55][117]=1;ram[55][118]=1;ram[55][119]=0;ram[55][120]=1;ram[55][121]=1;ram[55][122]=1;ram[55][123]=1;ram[55][124]=1;ram[55][125]=1;ram[55][126]=1;ram[55][127]=1;ram[55][128]=1;ram[55][129]=1;ram[55][130]=1;ram[55][131]=1;ram[55][132]=1;ram[55][133]=0;ram[55][134]=1;ram[55][135]=1;ram[55][136]=1;
        ram[56][0]=1;ram[56][1]=1;ram[56][2]=0;ram[56][3]=0;ram[56][4]=1;ram[56][5]=0;ram[56][6]=1;ram[56][7]=1;ram[56][8]=1;ram[56][9]=1;ram[56][10]=1;ram[56][11]=1;ram[56][12]=1;ram[56][13]=0;ram[56][14]=0;ram[56][15]=1;ram[56][16]=1;ram[56][17]=1;ram[56][18]=1;ram[56][19]=1;ram[56][20]=0;ram[56][21]=1;ram[56][22]=0;ram[56][23]=1;ram[56][24]=1;ram[56][25]=1;ram[56][26]=0;ram[56][27]=0;ram[56][28]=0;ram[56][29]=1;ram[56][30]=1;ram[56][31]=1;ram[56][32]=0;ram[56][33]=1;ram[56][34]=1;ram[56][35]=0;ram[56][36]=1;ram[56][37]=1;ram[56][38]=1;ram[56][39]=1;ram[56][40]=1;ram[56][41]=0;ram[56][42]=0;ram[56][43]=1;ram[56][44]=1;ram[56][45]=1;ram[56][46]=1;ram[56][47]=1;ram[56][48]=1;ram[56][49]=0;ram[56][50]=1;ram[56][51]=1;ram[56][52]=1;ram[56][53]=1;ram[56][54]=1;ram[56][55]=1;ram[56][56]=1;ram[56][57]=1;ram[56][58]=1;ram[56][59]=1;ram[56][60]=1;ram[56][61]=1;ram[56][62]=0;ram[56][63]=1;ram[56][64]=1;ram[56][65]=0;ram[56][66]=1;ram[56][67]=0;ram[56][68]=0;ram[56][69]=1;ram[56][70]=1;ram[56][71]=1;ram[56][72]=0;ram[56][73]=1;ram[56][74]=1;ram[56][75]=0;ram[56][76]=0;ram[56][77]=0;ram[56][78]=0;ram[56][79]=0;ram[56][80]=0;ram[56][81]=1;ram[56][82]=1;ram[56][83]=1;ram[56][84]=0;ram[56][85]=1;ram[56][86]=1;ram[56][87]=1;ram[56][88]=0;ram[56][89]=0;ram[56][90]=1;ram[56][91]=0;ram[56][92]=0;ram[56][93]=0;ram[56][94]=0;ram[56][95]=1;ram[56][96]=1;ram[56][97]=0;ram[56][98]=1;ram[56][99]=1;ram[56][100]=1;ram[56][101]=1;ram[56][102]=0;ram[56][103]=0;ram[56][104]=0;ram[56][105]=1;ram[56][106]=1;ram[56][107]=1;ram[56][108]=1;ram[56][109]=1;ram[56][110]=1;ram[56][111]=1;ram[56][112]=0;ram[56][113]=1;ram[56][114]=1;ram[56][115]=1;ram[56][116]=1;ram[56][117]=1;ram[56][118]=1;ram[56][119]=1;ram[56][120]=1;ram[56][121]=0;ram[56][122]=0;ram[56][123]=1;ram[56][124]=1;ram[56][125]=1;ram[56][126]=1;ram[56][127]=0;ram[56][128]=1;ram[56][129]=1;ram[56][130]=1;ram[56][131]=0;ram[56][132]=1;ram[56][133]=0;ram[56][134]=1;ram[56][135]=0;ram[56][136]=1;
        ram[57][0]=1;ram[57][1]=1;ram[57][2]=1;ram[57][3]=1;ram[57][4]=1;ram[57][5]=1;ram[57][6]=1;ram[57][7]=1;ram[57][8]=0;ram[57][9]=1;ram[57][10]=0;ram[57][11]=1;ram[57][12]=0;ram[57][13]=1;ram[57][14]=1;ram[57][15]=1;ram[57][16]=0;ram[57][17]=0;ram[57][18]=1;ram[57][19]=1;ram[57][20]=1;ram[57][21]=0;ram[57][22]=1;ram[57][23]=1;ram[57][24]=1;ram[57][25]=0;ram[57][26]=1;ram[57][27]=1;ram[57][28]=1;ram[57][29]=1;ram[57][30]=1;ram[57][31]=1;ram[57][32]=1;ram[57][33]=1;ram[57][34]=0;ram[57][35]=1;ram[57][36]=0;ram[57][37]=0;ram[57][38]=0;ram[57][39]=1;ram[57][40]=1;ram[57][41]=1;ram[57][42]=1;ram[57][43]=0;ram[57][44]=1;ram[57][45]=1;ram[57][46]=1;ram[57][47]=1;ram[57][48]=0;ram[57][49]=1;ram[57][50]=1;ram[57][51]=0;ram[57][52]=0;ram[57][53]=0;ram[57][54]=1;ram[57][55]=1;ram[57][56]=0;ram[57][57]=1;ram[57][58]=0;ram[57][59]=0;ram[57][60]=1;ram[57][61]=0;ram[57][62]=1;ram[57][63]=1;ram[57][64]=0;ram[57][65]=1;ram[57][66]=0;ram[57][67]=0;ram[57][68]=0;ram[57][69]=0;ram[57][70]=0;ram[57][71]=1;ram[57][72]=1;ram[57][73]=1;ram[57][74]=0;ram[57][75]=1;ram[57][76]=0;ram[57][77]=1;ram[57][78]=1;ram[57][79]=1;ram[57][80]=1;ram[57][81]=1;ram[57][82]=1;ram[57][83]=1;ram[57][84]=1;ram[57][85]=1;ram[57][86]=1;ram[57][87]=1;ram[57][88]=1;ram[57][89]=1;ram[57][90]=0;ram[57][91]=1;ram[57][92]=0;ram[57][93]=1;ram[57][94]=1;ram[57][95]=1;ram[57][96]=1;ram[57][97]=0;ram[57][98]=0;ram[57][99]=1;ram[57][100]=0;ram[57][101]=0;ram[57][102]=0;ram[57][103]=1;ram[57][104]=0;ram[57][105]=1;ram[57][106]=0;ram[57][107]=1;ram[57][108]=0;ram[57][109]=1;ram[57][110]=1;ram[57][111]=1;ram[57][112]=0;ram[57][113]=1;ram[57][114]=1;ram[57][115]=0;ram[57][116]=1;ram[57][117]=0;ram[57][118]=0;ram[57][119]=1;ram[57][120]=1;ram[57][121]=0;ram[57][122]=1;ram[57][123]=1;ram[57][124]=1;ram[57][125]=1;ram[57][126]=1;ram[57][127]=0;ram[57][128]=0;ram[57][129]=1;ram[57][130]=0;ram[57][131]=1;ram[57][132]=1;ram[57][133]=1;ram[57][134]=1;ram[57][135]=0;ram[57][136]=0;
        ram[58][0]=1;ram[58][1]=0;ram[58][2]=1;ram[58][3]=0;ram[58][4]=1;ram[58][5]=0;ram[58][6]=0;ram[58][7]=1;ram[58][8]=1;ram[58][9]=1;ram[58][10]=0;ram[58][11]=1;ram[58][12]=1;ram[58][13]=1;ram[58][14]=1;ram[58][15]=1;ram[58][16]=0;ram[58][17]=1;ram[58][18]=0;ram[58][19]=0;ram[58][20]=0;ram[58][21]=1;ram[58][22]=1;ram[58][23]=1;ram[58][24]=1;ram[58][25]=1;ram[58][26]=0;ram[58][27]=1;ram[58][28]=1;ram[58][29]=1;ram[58][30]=1;ram[58][31]=1;ram[58][32]=0;ram[58][33]=1;ram[58][34]=0;ram[58][35]=1;ram[58][36]=1;ram[58][37]=1;ram[58][38]=0;ram[58][39]=1;ram[58][40]=0;ram[58][41]=0;ram[58][42]=1;ram[58][43]=1;ram[58][44]=0;ram[58][45]=1;ram[58][46]=1;ram[58][47]=1;ram[58][48]=0;ram[58][49]=0;ram[58][50]=1;ram[58][51]=0;ram[58][52]=1;ram[58][53]=0;ram[58][54]=1;ram[58][55]=1;ram[58][56]=0;ram[58][57]=1;ram[58][58]=0;ram[58][59]=1;ram[58][60]=0;ram[58][61]=1;ram[58][62]=1;ram[58][63]=0;ram[58][64]=0;ram[58][65]=1;ram[58][66]=1;ram[58][67]=1;ram[58][68]=0;ram[58][69]=1;ram[58][70]=1;ram[58][71]=1;ram[58][72]=1;ram[58][73]=1;ram[58][74]=0;ram[58][75]=0;ram[58][76]=0;ram[58][77]=1;ram[58][78]=1;ram[58][79]=1;ram[58][80]=1;ram[58][81]=1;ram[58][82]=1;ram[58][83]=1;ram[58][84]=0;ram[58][85]=1;ram[58][86]=0;ram[58][87]=1;ram[58][88]=1;ram[58][89]=0;ram[58][90]=1;ram[58][91]=1;ram[58][92]=0;ram[58][93]=0;ram[58][94]=1;ram[58][95]=0;ram[58][96]=0;ram[58][97]=1;ram[58][98]=1;ram[58][99]=0;ram[58][100]=0;ram[58][101]=0;ram[58][102]=1;ram[58][103]=0;ram[58][104]=0;ram[58][105]=0;ram[58][106]=0;ram[58][107]=0;ram[58][108]=0;ram[58][109]=0;ram[58][110]=1;ram[58][111]=1;ram[58][112]=1;ram[58][113]=0;ram[58][114]=1;ram[58][115]=1;ram[58][116]=0;ram[58][117]=1;ram[58][118]=0;ram[58][119]=1;ram[58][120]=1;ram[58][121]=1;ram[58][122]=1;ram[58][123]=0;ram[58][124]=0;ram[58][125]=0;ram[58][126]=0;ram[58][127]=1;ram[58][128]=0;ram[58][129]=1;ram[58][130]=0;ram[58][131]=1;ram[58][132]=0;ram[58][133]=0;ram[58][134]=1;ram[58][135]=1;ram[58][136]=1;
        ram[59][0]=1;ram[59][1]=0;ram[59][2]=1;ram[59][3]=0;ram[59][4]=1;ram[59][5]=1;ram[59][6]=0;ram[59][7]=0;ram[59][8]=0;ram[59][9]=1;ram[59][10]=1;ram[59][11]=1;ram[59][12]=1;ram[59][13]=1;ram[59][14]=1;ram[59][15]=1;ram[59][16]=1;ram[59][17]=0;ram[59][18]=1;ram[59][19]=1;ram[59][20]=1;ram[59][21]=1;ram[59][22]=0;ram[59][23]=1;ram[59][24]=1;ram[59][25]=0;ram[59][26]=1;ram[59][27]=1;ram[59][28]=0;ram[59][29]=1;ram[59][30]=1;ram[59][31]=1;ram[59][32]=1;ram[59][33]=1;ram[59][34]=0;ram[59][35]=0;ram[59][36]=0;ram[59][37]=1;ram[59][38]=1;ram[59][39]=0;ram[59][40]=1;ram[59][41]=0;ram[59][42]=1;ram[59][43]=1;ram[59][44]=1;ram[59][45]=0;ram[59][46]=1;ram[59][47]=1;ram[59][48]=0;ram[59][49]=0;ram[59][50]=0;ram[59][51]=1;ram[59][52]=1;ram[59][53]=0;ram[59][54]=1;ram[59][55]=0;ram[59][56]=0;ram[59][57]=1;ram[59][58]=0;ram[59][59]=1;ram[59][60]=1;ram[59][61]=1;ram[59][62]=0;ram[59][63]=1;ram[59][64]=0;ram[59][65]=1;ram[59][66]=0;ram[59][67]=1;ram[59][68]=1;ram[59][69]=0;ram[59][70]=1;ram[59][71]=1;ram[59][72]=0;ram[59][73]=0;ram[59][74]=1;ram[59][75]=0;ram[59][76]=1;ram[59][77]=1;ram[59][78]=0;ram[59][79]=1;ram[59][80]=0;ram[59][81]=0;ram[59][82]=1;ram[59][83]=1;ram[59][84]=0;ram[59][85]=1;ram[59][86]=1;ram[59][87]=1;ram[59][88]=1;ram[59][89]=0;ram[59][90]=1;ram[59][91]=0;ram[59][92]=0;ram[59][93]=0;ram[59][94]=1;ram[59][95]=1;ram[59][96]=1;ram[59][97]=1;ram[59][98]=1;ram[59][99]=1;ram[59][100]=0;ram[59][101]=0;ram[59][102]=1;ram[59][103]=1;ram[59][104]=0;ram[59][105]=0;ram[59][106]=1;ram[59][107]=0;ram[59][108]=1;ram[59][109]=0;ram[59][110]=0;ram[59][111]=1;ram[59][112]=0;ram[59][113]=0;ram[59][114]=1;ram[59][115]=1;ram[59][116]=0;ram[59][117]=1;ram[59][118]=0;ram[59][119]=1;ram[59][120]=1;ram[59][121]=1;ram[59][122]=1;ram[59][123]=0;ram[59][124]=1;ram[59][125]=0;ram[59][126]=0;ram[59][127]=1;ram[59][128]=1;ram[59][129]=0;ram[59][130]=1;ram[59][131]=0;ram[59][132]=0;ram[59][133]=0;ram[59][134]=0;ram[59][135]=1;ram[59][136]=0;
        ram[60][0]=0;ram[60][1]=1;ram[60][2]=0;ram[60][3]=0;ram[60][4]=1;ram[60][5]=1;ram[60][6]=1;ram[60][7]=1;ram[60][8]=1;ram[60][9]=0;ram[60][10]=0;ram[60][11]=1;ram[60][12]=1;ram[60][13]=1;ram[60][14]=1;ram[60][15]=0;ram[60][16]=0;ram[60][17]=1;ram[60][18]=1;ram[60][19]=1;ram[60][20]=1;ram[60][21]=1;ram[60][22]=0;ram[60][23]=1;ram[60][24]=1;ram[60][25]=1;ram[60][26]=1;ram[60][27]=0;ram[60][28]=1;ram[60][29]=1;ram[60][30]=1;ram[60][31]=1;ram[60][32]=0;ram[60][33]=1;ram[60][34]=1;ram[60][35]=0;ram[60][36]=1;ram[60][37]=1;ram[60][38]=0;ram[60][39]=0;ram[60][40]=1;ram[60][41]=1;ram[60][42]=1;ram[60][43]=0;ram[60][44]=1;ram[60][45]=1;ram[60][46]=1;ram[60][47]=1;ram[60][48]=0;ram[60][49]=0;ram[60][50]=0;ram[60][51]=0;ram[60][52]=0;ram[60][53]=0;ram[60][54]=1;ram[60][55]=1;ram[60][56]=1;ram[60][57]=1;ram[60][58]=1;ram[60][59]=1;ram[60][60]=1;ram[60][61]=1;ram[60][62]=1;ram[60][63]=1;ram[60][64]=1;ram[60][65]=1;ram[60][66]=0;ram[60][67]=1;ram[60][68]=1;ram[60][69]=0;ram[60][70]=0;ram[60][71]=0;ram[60][72]=0;ram[60][73]=1;ram[60][74]=1;ram[60][75]=1;ram[60][76]=0;ram[60][77]=1;ram[60][78]=0;ram[60][79]=1;ram[60][80]=1;ram[60][81]=1;ram[60][82]=1;ram[60][83]=0;ram[60][84]=1;ram[60][85]=1;ram[60][86]=0;ram[60][87]=0;ram[60][88]=0;ram[60][89]=1;ram[60][90]=1;ram[60][91]=0;ram[60][92]=0;ram[60][93]=1;ram[60][94]=1;ram[60][95]=1;ram[60][96]=1;ram[60][97]=0;ram[60][98]=0;ram[60][99]=0;ram[60][100]=1;ram[60][101]=1;ram[60][102]=0;ram[60][103]=1;ram[60][104]=1;ram[60][105]=1;ram[60][106]=1;ram[60][107]=0;ram[60][108]=1;ram[60][109]=1;ram[60][110]=0;ram[60][111]=1;ram[60][112]=1;ram[60][113]=1;ram[60][114]=1;ram[60][115]=1;ram[60][116]=0;ram[60][117]=0;ram[60][118]=1;ram[60][119]=1;ram[60][120]=1;ram[60][121]=1;ram[60][122]=0;ram[60][123]=0;ram[60][124]=1;ram[60][125]=0;ram[60][126]=1;ram[60][127]=0;ram[60][128]=1;ram[60][129]=0;ram[60][130]=1;ram[60][131]=1;ram[60][132]=0;ram[60][133]=0;ram[60][134]=0;ram[60][135]=0;ram[60][136]=1;
        ram[61][0]=1;ram[61][1]=0;ram[61][2]=1;ram[61][3]=0;ram[61][4]=1;ram[61][5]=0;ram[61][6]=1;ram[61][7]=1;ram[61][8]=0;ram[61][9]=1;ram[61][10]=1;ram[61][11]=0;ram[61][12]=0;ram[61][13]=1;ram[61][14]=1;ram[61][15]=0;ram[61][16]=1;ram[61][17]=0;ram[61][18]=1;ram[61][19]=1;ram[61][20]=1;ram[61][21]=1;ram[61][22]=1;ram[61][23]=1;ram[61][24]=1;ram[61][25]=1;ram[61][26]=1;ram[61][27]=0;ram[61][28]=1;ram[61][29]=1;ram[61][30]=1;ram[61][31]=1;ram[61][32]=1;ram[61][33]=1;ram[61][34]=1;ram[61][35]=0;ram[61][36]=1;ram[61][37]=1;ram[61][38]=1;ram[61][39]=1;ram[61][40]=0;ram[61][41]=0;ram[61][42]=1;ram[61][43]=1;ram[61][44]=0;ram[61][45]=1;ram[61][46]=0;ram[61][47]=1;ram[61][48]=0;ram[61][49]=0;ram[61][50]=1;ram[61][51]=1;ram[61][52]=1;ram[61][53]=0;ram[61][54]=0;ram[61][55]=1;ram[61][56]=1;ram[61][57]=1;ram[61][58]=1;ram[61][59]=1;ram[61][60]=1;ram[61][61]=1;ram[61][62]=1;ram[61][63]=1;ram[61][64]=0;ram[61][65]=1;ram[61][66]=0;ram[61][67]=1;ram[61][68]=1;ram[61][69]=1;ram[61][70]=0;ram[61][71]=1;ram[61][72]=0;ram[61][73]=0;ram[61][74]=1;ram[61][75]=1;ram[61][76]=0;ram[61][77]=1;ram[61][78]=1;ram[61][79]=0;ram[61][80]=1;ram[61][81]=1;ram[61][82]=0;ram[61][83]=1;ram[61][84]=1;ram[61][85]=0;ram[61][86]=1;ram[61][87]=0;ram[61][88]=1;ram[61][89]=0;ram[61][90]=1;ram[61][91]=1;ram[61][92]=1;ram[61][93]=1;ram[61][94]=1;ram[61][95]=0;ram[61][96]=1;ram[61][97]=0;ram[61][98]=1;ram[61][99]=1;ram[61][100]=1;ram[61][101]=1;ram[61][102]=0;ram[61][103]=0;ram[61][104]=1;ram[61][105]=1;ram[61][106]=0;ram[61][107]=1;ram[61][108]=0;ram[61][109]=1;ram[61][110]=1;ram[61][111]=0;ram[61][112]=0;ram[61][113]=1;ram[61][114]=1;ram[61][115]=0;ram[61][116]=1;ram[61][117]=0;ram[61][118]=1;ram[61][119]=0;ram[61][120]=0;ram[61][121]=0;ram[61][122]=0;ram[61][123]=1;ram[61][124]=0;ram[61][125]=0;ram[61][126]=0;ram[61][127]=1;ram[61][128]=1;ram[61][129]=0;ram[61][130]=1;ram[61][131]=1;ram[61][132]=1;ram[61][133]=0;ram[61][134]=1;ram[61][135]=1;ram[61][136]=0;
        ram[62][0]=1;ram[62][1]=1;ram[62][2]=1;ram[62][3]=1;ram[62][4]=0;ram[62][5]=1;ram[62][6]=1;ram[62][7]=1;ram[62][8]=0;ram[62][9]=0;ram[62][10]=1;ram[62][11]=0;ram[62][12]=1;ram[62][13]=0;ram[62][14]=1;ram[62][15]=1;ram[62][16]=1;ram[62][17]=0;ram[62][18]=1;ram[62][19]=0;ram[62][20]=1;ram[62][21]=1;ram[62][22]=1;ram[62][23]=1;ram[62][24]=1;ram[62][25]=1;ram[62][26]=1;ram[62][27]=1;ram[62][28]=1;ram[62][29]=1;ram[62][30]=1;ram[62][31]=1;ram[62][32]=1;ram[62][33]=1;ram[62][34]=1;ram[62][35]=0;ram[62][36]=1;ram[62][37]=1;ram[62][38]=0;ram[62][39]=1;ram[62][40]=1;ram[62][41]=1;ram[62][42]=0;ram[62][43]=1;ram[62][44]=1;ram[62][45]=0;ram[62][46]=1;ram[62][47]=1;ram[62][48]=1;ram[62][49]=1;ram[62][50]=1;ram[62][51]=1;ram[62][52]=1;ram[62][53]=0;ram[62][54]=0;ram[62][55]=0;ram[62][56]=0;ram[62][57]=0;ram[62][58]=1;ram[62][59]=1;ram[62][60]=0;ram[62][61]=1;ram[62][62]=1;ram[62][63]=1;ram[62][64]=1;ram[62][65]=1;ram[62][66]=1;ram[62][67]=1;ram[62][68]=1;ram[62][69]=0;ram[62][70]=0;ram[62][71]=1;ram[62][72]=1;ram[62][73]=1;ram[62][74]=0;ram[62][75]=1;ram[62][76]=0;ram[62][77]=1;ram[62][78]=0;ram[62][79]=1;ram[62][80]=1;ram[62][81]=1;ram[62][82]=1;ram[62][83]=0;ram[62][84]=1;ram[62][85]=1;ram[62][86]=0;ram[62][87]=1;ram[62][88]=1;ram[62][89]=1;ram[62][90]=1;ram[62][91]=1;ram[62][92]=0;ram[62][93]=1;ram[62][94]=1;ram[62][95]=0;ram[62][96]=1;ram[62][97]=0;ram[62][98]=1;ram[62][99]=0;ram[62][100]=0;ram[62][101]=1;ram[62][102]=1;ram[62][103]=1;ram[62][104]=1;ram[62][105]=0;ram[62][106]=1;ram[62][107]=1;ram[62][108]=0;ram[62][109]=1;ram[62][110]=1;ram[62][111]=0;ram[62][112]=1;ram[62][113]=1;ram[62][114]=1;ram[62][115]=1;ram[62][116]=1;ram[62][117]=1;ram[62][118]=1;ram[62][119]=1;ram[62][120]=1;ram[62][121]=0;ram[62][122]=1;ram[62][123]=1;ram[62][124]=0;ram[62][125]=0;ram[62][126]=1;ram[62][127]=0;ram[62][128]=1;ram[62][129]=1;ram[62][130]=1;ram[62][131]=0;ram[62][132]=0;ram[62][133]=0;ram[62][134]=1;ram[62][135]=1;ram[62][136]=1;
        ram[63][0]=1;ram[63][1]=1;ram[63][2]=0;ram[63][3]=1;ram[63][4]=0;ram[63][5]=0;ram[63][6]=1;ram[63][7]=1;ram[63][8]=1;ram[63][9]=1;ram[63][10]=0;ram[63][11]=0;ram[63][12]=0;ram[63][13]=1;ram[63][14]=0;ram[63][15]=1;ram[63][16]=0;ram[63][17]=1;ram[63][18]=0;ram[63][19]=0;ram[63][20]=1;ram[63][21]=1;ram[63][22]=1;ram[63][23]=1;ram[63][24]=1;ram[63][25]=1;ram[63][26]=0;ram[63][27]=0;ram[63][28]=1;ram[63][29]=1;ram[63][30]=1;ram[63][31]=1;ram[63][32]=0;ram[63][33]=0;ram[63][34]=1;ram[63][35]=0;ram[63][36]=1;ram[63][37]=1;ram[63][38]=0;ram[63][39]=1;ram[63][40]=0;ram[63][41]=0;ram[63][42]=1;ram[63][43]=1;ram[63][44]=1;ram[63][45]=0;ram[63][46]=0;ram[63][47]=1;ram[63][48]=1;ram[63][49]=1;ram[63][50]=1;ram[63][51]=1;ram[63][52]=0;ram[63][53]=0;ram[63][54]=1;ram[63][55]=0;ram[63][56]=1;ram[63][57]=0;ram[63][58]=0;ram[63][59]=1;ram[63][60]=1;ram[63][61]=1;ram[63][62]=1;ram[63][63]=0;ram[63][64]=1;ram[63][65]=1;ram[63][66]=1;ram[63][67]=0;ram[63][68]=0;ram[63][69]=1;ram[63][70]=0;ram[63][71]=0;ram[63][72]=1;ram[63][73]=0;ram[63][74]=0;ram[63][75]=1;ram[63][76]=0;ram[63][77]=1;ram[63][78]=1;ram[63][79]=1;ram[63][80]=1;ram[63][81]=0;ram[63][82]=0;ram[63][83]=1;ram[63][84]=1;ram[63][85]=0;ram[63][86]=1;ram[63][87]=1;ram[63][88]=1;ram[63][89]=1;ram[63][90]=0;ram[63][91]=1;ram[63][92]=0;ram[63][93]=1;ram[63][94]=1;ram[63][95]=1;ram[63][96]=1;ram[63][97]=0;ram[63][98]=0;ram[63][99]=1;ram[63][100]=0;ram[63][101]=0;ram[63][102]=1;ram[63][103]=1;ram[63][104]=0;ram[63][105]=1;ram[63][106]=1;ram[63][107]=1;ram[63][108]=1;ram[63][109]=0;ram[63][110]=1;ram[63][111]=1;ram[63][112]=0;ram[63][113]=0;ram[63][114]=1;ram[63][115]=1;ram[63][116]=0;ram[63][117]=0;ram[63][118]=1;ram[63][119]=1;ram[63][120]=0;ram[63][121]=0;ram[63][122]=0;ram[63][123]=0;ram[63][124]=0;ram[63][125]=1;ram[63][126]=1;ram[63][127]=1;ram[63][128]=1;ram[63][129]=1;ram[63][130]=0;ram[63][131]=0;ram[63][132]=0;ram[63][133]=0;ram[63][134]=1;ram[63][135]=1;ram[63][136]=0;
        ram[64][0]=1;ram[64][1]=1;ram[64][2]=1;ram[64][3]=1;ram[64][4]=1;ram[64][5]=1;ram[64][6]=1;ram[64][7]=1;ram[64][8]=0;ram[64][9]=0;ram[64][10]=0;ram[64][11]=0;ram[64][12]=0;ram[64][13]=1;ram[64][14]=1;ram[64][15]=0;ram[64][16]=1;ram[64][17]=0;ram[64][18]=1;ram[64][19]=0;ram[64][20]=1;ram[64][21]=1;ram[64][22]=0;ram[64][23]=0;ram[64][24]=1;ram[64][25]=1;ram[64][26]=1;ram[64][27]=0;ram[64][28]=0;ram[64][29]=0;ram[64][30]=0;ram[64][31]=0;ram[64][32]=1;ram[64][33]=1;ram[64][34]=1;ram[64][35]=1;ram[64][36]=1;ram[64][37]=1;ram[64][38]=1;ram[64][39]=1;ram[64][40]=0;ram[64][41]=1;ram[64][42]=1;ram[64][43]=1;ram[64][44]=0;ram[64][45]=1;ram[64][46]=1;ram[64][47]=1;ram[64][48]=1;ram[64][49]=0;ram[64][50]=1;ram[64][51]=1;ram[64][52]=1;ram[64][53]=1;ram[64][54]=0;ram[64][55]=1;ram[64][56]=1;ram[64][57]=0;ram[64][58]=1;ram[64][59]=1;ram[64][60]=0;ram[64][61]=1;ram[64][62]=1;ram[64][63]=1;ram[64][64]=0;ram[64][65]=0;ram[64][66]=1;ram[64][67]=1;ram[64][68]=1;ram[64][69]=0;ram[64][70]=0;ram[64][71]=0;ram[64][72]=1;ram[64][73]=1;ram[64][74]=0;ram[64][75]=1;ram[64][76]=0;ram[64][77]=1;ram[64][78]=0;ram[64][79]=1;ram[64][80]=1;ram[64][81]=1;ram[64][82]=0;ram[64][83]=1;ram[64][84]=1;ram[64][85]=1;ram[64][86]=0;ram[64][87]=1;ram[64][88]=0;ram[64][89]=0;ram[64][90]=1;ram[64][91]=0;ram[64][92]=1;ram[64][93]=0;ram[64][94]=1;ram[64][95]=1;ram[64][96]=1;ram[64][97]=0;ram[64][98]=0;ram[64][99]=1;ram[64][100]=1;ram[64][101]=0;ram[64][102]=0;ram[64][103]=1;ram[64][104]=1;ram[64][105]=1;ram[64][106]=0;ram[64][107]=1;ram[64][108]=0;ram[64][109]=1;ram[64][110]=1;ram[64][111]=1;ram[64][112]=1;ram[64][113]=0;ram[64][114]=0;ram[64][115]=0;ram[64][116]=1;ram[64][117]=1;ram[64][118]=0;ram[64][119]=0;ram[64][120]=0;ram[64][121]=0;ram[64][122]=1;ram[64][123]=1;ram[64][124]=1;ram[64][125]=1;ram[64][126]=1;ram[64][127]=1;ram[64][128]=0;ram[64][129]=0;ram[64][130]=1;ram[64][131]=1;ram[64][132]=0;ram[64][133]=0;ram[64][134]=1;ram[64][135]=1;ram[64][136]=0;
        ram[65][0]=0;ram[65][1]=1;ram[65][2]=0;ram[65][3]=1;ram[65][4]=1;ram[65][5]=0;ram[65][6]=1;ram[65][7]=1;ram[65][8]=1;ram[65][9]=0;ram[65][10]=0;ram[65][11]=1;ram[65][12]=1;ram[65][13]=1;ram[65][14]=0;ram[65][15]=0;ram[65][16]=1;ram[65][17]=0;ram[65][18]=1;ram[65][19]=0;ram[65][20]=0;ram[65][21]=0;ram[65][22]=1;ram[65][23]=1;ram[65][24]=1;ram[65][25]=1;ram[65][26]=1;ram[65][27]=1;ram[65][28]=0;ram[65][29]=1;ram[65][30]=0;ram[65][31]=0;ram[65][32]=0;ram[65][33]=1;ram[65][34]=1;ram[65][35]=1;ram[65][36]=1;ram[65][37]=0;ram[65][38]=1;ram[65][39]=1;ram[65][40]=1;ram[65][41]=1;ram[65][42]=1;ram[65][43]=1;ram[65][44]=0;ram[65][45]=0;ram[65][46]=1;ram[65][47]=1;ram[65][48]=1;ram[65][49]=0;ram[65][50]=1;ram[65][51]=0;ram[65][52]=1;ram[65][53]=1;ram[65][54]=0;ram[65][55]=1;ram[65][56]=0;ram[65][57]=0;ram[65][58]=0;ram[65][59]=1;ram[65][60]=1;ram[65][61]=0;ram[65][62]=0;ram[65][63]=1;ram[65][64]=1;ram[65][65]=1;ram[65][66]=0;ram[65][67]=1;ram[65][68]=1;ram[65][69]=0;ram[65][70]=1;ram[65][71]=1;ram[65][72]=1;ram[65][73]=0;ram[65][74]=0;ram[65][75]=0;ram[65][76]=1;ram[65][77]=0;ram[65][78]=0;ram[65][79]=1;ram[65][80]=1;ram[65][81]=0;ram[65][82]=1;ram[65][83]=1;ram[65][84]=1;ram[65][85]=0;ram[65][86]=0;ram[65][87]=1;ram[65][88]=1;ram[65][89]=1;ram[65][90]=0;ram[65][91]=1;ram[65][92]=0;ram[65][93]=1;ram[65][94]=1;ram[65][95]=0;ram[65][96]=1;ram[65][97]=1;ram[65][98]=1;ram[65][99]=1;ram[65][100]=1;ram[65][101]=0;ram[65][102]=1;ram[65][103]=1;ram[65][104]=1;ram[65][105]=1;ram[65][106]=1;ram[65][107]=0;ram[65][108]=0;ram[65][109]=1;ram[65][110]=0;ram[65][111]=1;ram[65][112]=0;ram[65][113]=1;ram[65][114]=0;ram[65][115]=1;ram[65][116]=1;ram[65][117]=0;ram[65][118]=0;ram[65][119]=0;ram[65][120]=0;ram[65][121]=0;ram[65][122]=0;ram[65][123]=1;ram[65][124]=0;ram[65][125]=1;ram[65][126]=0;ram[65][127]=1;ram[65][128]=0;ram[65][129]=1;ram[65][130]=1;ram[65][131]=0;ram[65][132]=0;ram[65][133]=1;ram[65][134]=1;ram[65][135]=1;ram[65][136]=1;
        ram[66][0]=1;ram[66][1]=1;ram[66][2]=1;ram[66][3]=1;ram[66][4]=1;ram[66][5]=1;ram[66][6]=0;ram[66][7]=1;ram[66][8]=1;ram[66][9]=1;ram[66][10]=0;ram[66][11]=1;ram[66][12]=0;ram[66][13]=0;ram[66][14]=1;ram[66][15]=1;ram[66][16]=1;ram[66][17]=1;ram[66][18]=1;ram[66][19]=1;ram[66][20]=0;ram[66][21]=1;ram[66][22]=1;ram[66][23]=1;ram[66][24]=1;ram[66][25]=0;ram[66][26]=1;ram[66][27]=1;ram[66][28]=1;ram[66][29]=1;ram[66][30]=1;ram[66][31]=0;ram[66][32]=1;ram[66][33]=0;ram[66][34]=1;ram[66][35]=0;ram[66][36]=1;ram[66][37]=0;ram[66][38]=0;ram[66][39]=1;ram[66][40]=1;ram[66][41]=0;ram[66][42]=1;ram[66][43]=0;ram[66][44]=0;ram[66][45]=0;ram[66][46]=1;ram[66][47]=0;ram[66][48]=1;ram[66][49]=1;ram[66][50]=1;ram[66][51]=1;ram[66][52]=1;ram[66][53]=1;ram[66][54]=1;ram[66][55]=1;ram[66][56]=1;ram[66][57]=1;ram[66][58]=0;ram[66][59]=1;ram[66][60]=1;ram[66][61]=1;ram[66][62]=1;ram[66][63]=0;ram[66][64]=0;ram[66][65]=0;ram[66][66]=0;ram[66][67]=1;ram[66][68]=1;ram[66][69]=1;ram[66][70]=1;ram[66][71]=1;ram[66][72]=1;ram[66][73]=1;ram[66][74]=1;ram[66][75]=1;ram[66][76]=0;ram[66][77]=1;ram[66][78]=1;ram[66][79]=0;ram[66][80]=1;ram[66][81]=1;ram[66][82]=0;ram[66][83]=0;ram[66][84]=0;ram[66][85]=0;ram[66][86]=1;ram[66][87]=0;ram[66][88]=1;ram[66][89]=0;ram[66][90]=1;ram[66][91]=1;ram[66][92]=0;ram[66][93]=1;ram[66][94]=1;ram[66][95]=1;ram[66][96]=1;ram[66][97]=0;ram[66][98]=1;ram[66][99]=0;ram[66][100]=1;ram[66][101]=0;ram[66][102]=1;ram[66][103]=1;ram[66][104]=0;ram[66][105]=1;ram[66][106]=1;ram[66][107]=1;ram[66][108]=1;ram[66][109]=1;ram[66][110]=0;ram[66][111]=0;ram[66][112]=0;ram[66][113]=0;ram[66][114]=1;ram[66][115]=0;ram[66][116]=0;ram[66][117]=1;ram[66][118]=0;ram[66][119]=0;ram[66][120]=1;ram[66][121]=1;ram[66][122]=1;ram[66][123]=1;ram[66][124]=1;ram[66][125]=0;ram[66][126]=1;ram[66][127]=1;ram[66][128]=1;ram[66][129]=1;ram[66][130]=1;ram[66][131]=1;ram[66][132]=1;ram[66][133]=0;ram[66][134]=1;ram[66][135]=1;ram[66][136]=0;
        ram[67][0]=1;ram[67][1]=1;ram[67][2]=0;ram[67][3]=1;ram[67][4]=1;ram[67][5]=1;ram[67][6]=0;ram[67][7]=0;ram[67][8]=1;ram[67][9]=1;ram[67][10]=0;ram[67][11]=1;ram[67][12]=1;ram[67][13]=0;ram[67][14]=1;ram[67][15]=1;ram[67][16]=1;ram[67][17]=0;ram[67][18]=0;ram[67][19]=0;ram[67][20]=1;ram[67][21]=0;ram[67][22]=0;ram[67][23]=0;ram[67][24]=0;ram[67][25]=0;ram[67][26]=1;ram[67][27]=1;ram[67][28]=1;ram[67][29]=1;ram[67][30]=1;ram[67][31]=1;ram[67][32]=1;ram[67][33]=1;ram[67][34]=1;ram[67][35]=0;ram[67][36]=1;ram[67][37]=1;ram[67][38]=0;ram[67][39]=1;ram[67][40]=1;ram[67][41]=0;ram[67][42]=1;ram[67][43]=0;ram[67][44]=1;ram[67][45]=1;ram[67][46]=1;ram[67][47]=1;ram[67][48]=1;ram[67][49]=1;ram[67][50]=1;ram[67][51]=1;ram[67][52]=1;ram[67][53]=0;ram[67][54]=1;ram[67][55]=0;ram[67][56]=1;ram[67][57]=1;ram[67][58]=0;ram[67][59]=1;ram[67][60]=1;ram[67][61]=0;ram[67][62]=0;ram[67][63]=1;ram[67][64]=0;ram[67][65]=0;ram[67][66]=0;ram[67][67]=1;ram[67][68]=1;ram[67][69]=0;ram[67][70]=1;ram[67][71]=0;ram[67][72]=1;ram[67][73]=1;ram[67][74]=1;ram[67][75]=1;ram[67][76]=1;ram[67][77]=1;ram[67][78]=1;ram[67][79]=0;ram[67][80]=1;ram[67][81]=1;ram[67][82]=1;ram[67][83]=1;ram[67][84]=1;ram[67][85]=0;ram[67][86]=1;ram[67][87]=1;ram[67][88]=1;ram[67][89]=0;ram[67][90]=0;ram[67][91]=0;ram[67][92]=1;ram[67][93]=1;ram[67][94]=0;ram[67][95]=1;ram[67][96]=1;ram[67][97]=0;ram[67][98]=1;ram[67][99]=1;ram[67][100]=1;ram[67][101]=1;ram[67][102]=1;ram[67][103]=1;ram[67][104]=1;ram[67][105]=0;ram[67][106]=1;ram[67][107]=1;ram[67][108]=0;ram[67][109]=1;ram[67][110]=0;ram[67][111]=1;ram[67][112]=0;ram[67][113]=1;ram[67][114]=1;ram[67][115]=1;ram[67][116]=1;ram[67][117]=1;ram[67][118]=0;ram[67][119]=1;ram[67][120]=1;ram[67][121]=0;ram[67][122]=0;ram[67][123]=1;ram[67][124]=1;ram[67][125]=1;ram[67][126]=1;ram[67][127]=0;ram[67][128]=1;ram[67][129]=0;ram[67][130]=1;ram[67][131]=0;ram[67][132]=1;ram[67][133]=1;ram[67][134]=1;ram[67][135]=0;ram[67][136]=1;
        ram[68][0]=1;ram[68][1]=1;ram[68][2]=1;ram[68][3]=1;ram[68][4]=1;ram[68][5]=1;ram[68][6]=1;ram[68][7]=0;ram[68][8]=1;ram[68][9]=0;ram[68][10]=1;ram[68][11]=1;ram[68][12]=1;ram[68][13]=0;ram[68][14]=1;ram[68][15]=0;ram[68][16]=1;ram[68][17]=0;ram[68][18]=1;ram[68][19]=1;ram[68][20]=1;ram[68][21]=1;ram[68][22]=0;ram[68][23]=1;ram[68][24]=0;ram[68][25]=0;ram[68][26]=1;ram[68][27]=1;ram[68][28]=1;ram[68][29]=0;ram[68][30]=0;ram[68][31]=0;ram[68][32]=0;ram[68][33]=1;ram[68][34]=0;ram[68][35]=0;ram[68][36]=0;ram[68][37]=0;ram[68][38]=0;ram[68][39]=0;ram[68][40]=0;ram[68][41]=0;ram[68][42]=0;ram[68][43]=0;ram[68][44]=1;ram[68][45]=0;ram[68][46]=1;ram[68][47]=0;ram[68][48]=0;ram[68][49]=1;ram[68][50]=1;ram[68][51]=0;ram[68][52]=1;ram[68][53]=0;ram[68][54]=1;ram[68][55]=1;ram[68][56]=1;ram[68][57]=1;ram[68][58]=0;ram[68][59]=1;ram[68][60]=0;ram[68][61]=1;ram[68][62]=1;ram[68][63]=1;ram[68][64]=0;ram[68][65]=0;ram[68][66]=0;ram[68][67]=1;ram[68][68]=0;ram[68][69]=0;ram[68][70]=0;ram[68][71]=1;ram[68][72]=0;ram[68][73]=0;ram[68][74]=0;ram[68][75]=0;ram[68][76]=1;ram[68][77]=0;ram[68][78]=0;ram[68][79]=1;ram[68][80]=0;ram[68][81]=0;ram[68][82]=1;ram[68][83]=0;ram[68][84]=0;ram[68][85]=1;ram[68][86]=1;ram[68][87]=0;ram[68][88]=1;ram[68][89]=1;ram[68][90]=1;ram[68][91]=0;ram[68][92]=1;ram[68][93]=1;ram[68][94]=0;ram[68][95]=1;ram[68][96]=1;ram[68][97]=0;ram[68][98]=1;ram[68][99]=0;ram[68][100]=0;ram[68][101]=0;ram[68][102]=1;ram[68][103]=1;ram[68][104]=1;ram[68][105]=0;ram[68][106]=1;ram[68][107]=0;ram[68][108]=1;ram[68][109]=1;ram[68][110]=1;ram[68][111]=1;ram[68][112]=1;ram[68][113]=0;ram[68][114]=1;ram[68][115]=1;ram[68][116]=1;ram[68][117]=0;ram[68][118]=1;ram[68][119]=1;ram[68][120]=0;ram[68][121]=1;ram[68][122]=0;ram[68][123]=1;ram[68][124]=0;ram[68][125]=0;ram[68][126]=0;ram[68][127]=0;ram[68][128]=1;ram[68][129]=1;ram[68][130]=1;ram[68][131]=1;ram[68][132]=1;ram[68][133]=0;ram[68][134]=1;ram[68][135]=1;ram[68][136]=1;
        ram[69][0]=1;ram[69][1]=1;ram[69][2]=1;ram[69][3]=1;ram[69][4]=0;ram[69][5]=0;ram[69][6]=1;ram[69][7]=1;ram[69][8]=1;ram[69][9]=1;ram[69][10]=1;ram[69][11]=0;ram[69][12]=1;ram[69][13]=0;ram[69][14]=0;ram[69][15]=1;ram[69][16]=1;ram[69][17]=1;ram[69][18]=1;ram[69][19]=0;ram[69][20]=1;ram[69][21]=0;ram[69][22]=1;ram[69][23]=0;ram[69][24]=0;ram[69][25]=1;ram[69][26]=0;ram[69][27]=0;ram[69][28]=1;ram[69][29]=1;ram[69][30]=1;ram[69][31]=1;ram[69][32]=1;ram[69][33]=1;ram[69][34]=0;ram[69][35]=1;ram[69][36]=0;ram[69][37]=1;ram[69][38]=1;ram[69][39]=1;ram[69][40]=1;ram[69][41]=1;ram[69][42]=1;ram[69][43]=1;ram[69][44]=1;ram[69][45]=1;ram[69][46]=0;ram[69][47]=1;ram[69][48]=1;ram[69][49]=1;ram[69][50]=1;ram[69][51]=1;ram[69][52]=0;ram[69][53]=1;ram[69][54]=1;ram[69][55]=0;ram[69][56]=0;ram[69][57]=1;ram[69][58]=1;ram[69][59]=1;ram[69][60]=1;ram[69][61]=0;ram[69][62]=1;ram[69][63]=1;ram[69][64]=0;ram[69][65]=0;ram[69][66]=1;ram[69][67]=1;ram[69][68]=1;ram[69][69]=1;ram[69][70]=1;ram[69][71]=1;ram[69][72]=0;ram[69][73]=1;ram[69][74]=1;ram[69][75]=1;ram[69][76]=0;ram[69][77]=0;ram[69][78]=0;ram[69][79]=1;ram[69][80]=1;ram[69][81]=1;ram[69][82]=1;ram[69][83]=1;ram[69][84]=1;ram[69][85]=0;ram[69][86]=1;ram[69][87]=0;ram[69][88]=1;ram[69][89]=0;ram[69][90]=1;ram[69][91]=1;ram[69][92]=1;ram[69][93]=1;ram[69][94]=1;ram[69][95]=0;ram[69][96]=1;ram[69][97]=1;ram[69][98]=1;ram[69][99]=1;ram[69][100]=1;ram[69][101]=1;ram[69][102]=1;ram[69][103]=1;ram[69][104]=1;ram[69][105]=1;ram[69][106]=1;ram[69][107]=0;ram[69][108]=0;ram[69][109]=1;ram[69][110]=1;ram[69][111]=0;ram[69][112]=0;ram[69][113]=1;ram[69][114]=0;ram[69][115]=0;ram[69][116]=1;ram[69][117]=1;ram[69][118]=0;ram[69][119]=0;ram[69][120]=0;ram[69][121]=1;ram[69][122]=1;ram[69][123]=0;ram[69][124]=0;ram[69][125]=0;ram[69][126]=0;ram[69][127]=1;ram[69][128]=1;ram[69][129]=0;ram[69][130]=1;ram[69][131]=0;ram[69][132]=1;ram[69][133]=1;ram[69][134]=1;ram[69][135]=0;ram[69][136]=0;
        ram[70][0]=1;ram[70][1]=1;ram[70][2]=0;ram[70][3]=1;ram[70][4]=1;ram[70][5]=1;ram[70][6]=0;ram[70][7]=0;ram[70][8]=0;ram[70][9]=0;ram[70][10]=1;ram[70][11]=0;ram[70][12]=1;ram[70][13]=1;ram[70][14]=0;ram[70][15]=1;ram[70][16]=1;ram[70][17]=0;ram[70][18]=1;ram[70][19]=1;ram[70][20]=0;ram[70][21]=0;ram[70][22]=1;ram[70][23]=0;ram[70][24]=0;ram[70][25]=0;ram[70][26]=0;ram[70][27]=0;ram[70][28]=0;ram[70][29]=1;ram[70][30]=0;ram[70][31]=1;ram[70][32]=1;ram[70][33]=1;ram[70][34]=1;ram[70][35]=1;ram[70][36]=1;ram[70][37]=1;ram[70][38]=0;ram[70][39]=0;ram[70][40]=1;ram[70][41]=1;ram[70][42]=1;ram[70][43]=1;ram[70][44]=1;ram[70][45]=1;ram[70][46]=1;ram[70][47]=1;ram[70][48]=1;ram[70][49]=1;ram[70][50]=1;ram[70][51]=1;ram[70][52]=0;ram[70][53]=1;ram[70][54]=0;ram[70][55]=0;ram[70][56]=1;ram[70][57]=1;ram[70][58]=1;ram[70][59]=1;ram[70][60]=1;ram[70][61]=1;ram[70][62]=1;ram[70][63]=0;ram[70][64]=0;ram[70][65]=1;ram[70][66]=1;ram[70][67]=1;ram[70][68]=1;ram[70][69]=1;ram[70][70]=0;ram[70][71]=0;ram[70][72]=1;ram[70][73]=1;ram[70][74]=1;ram[70][75]=1;ram[70][76]=0;ram[70][77]=1;ram[70][78]=1;ram[70][79]=1;ram[70][80]=0;ram[70][81]=0;ram[70][82]=1;ram[70][83]=1;ram[70][84]=1;ram[70][85]=1;ram[70][86]=1;ram[70][87]=0;ram[70][88]=1;ram[70][89]=0;ram[70][90]=0;ram[70][91]=1;ram[70][92]=1;ram[70][93]=0;ram[70][94]=1;ram[70][95]=1;ram[70][96]=1;ram[70][97]=1;ram[70][98]=1;ram[70][99]=1;ram[70][100]=1;ram[70][101]=1;ram[70][102]=1;ram[70][103]=1;ram[70][104]=1;ram[70][105]=0;ram[70][106]=1;ram[70][107]=0;ram[70][108]=1;ram[70][109]=1;ram[70][110]=1;ram[70][111]=1;ram[70][112]=1;ram[70][113]=0;ram[70][114]=1;ram[70][115]=1;ram[70][116]=1;ram[70][117]=0;ram[70][118]=1;ram[70][119]=0;ram[70][120]=1;ram[70][121]=0;ram[70][122]=0;ram[70][123]=1;ram[70][124]=0;ram[70][125]=1;ram[70][126]=1;ram[70][127]=1;ram[70][128]=0;ram[70][129]=0;ram[70][130]=1;ram[70][131]=1;ram[70][132]=0;ram[70][133]=1;ram[70][134]=1;ram[70][135]=0;ram[70][136]=1;
        ram[71][0]=1;ram[71][1]=1;ram[71][2]=1;ram[71][3]=0;ram[71][4]=0;ram[71][5]=1;ram[71][6]=1;ram[71][7]=0;ram[71][8]=1;ram[71][9]=0;ram[71][10]=1;ram[71][11]=1;ram[71][12]=0;ram[71][13]=0;ram[71][14]=1;ram[71][15]=1;ram[71][16]=0;ram[71][17]=0;ram[71][18]=1;ram[71][19]=0;ram[71][20]=0;ram[71][21]=1;ram[71][22]=1;ram[71][23]=1;ram[71][24]=1;ram[71][25]=1;ram[71][26]=1;ram[71][27]=0;ram[71][28]=0;ram[71][29]=1;ram[71][30]=0;ram[71][31]=0;ram[71][32]=1;ram[71][33]=1;ram[71][34]=0;ram[71][35]=1;ram[71][36]=1;ram[71][37]=1;ram[71][38]=1;ram[71][39]=1;ram[71][40]=0;ram[71][41]=1;ram[71][42]=0;ram[71][43]=0;ram[71][44]=1;ram[71][45]=0;ram[71][46]=1;ram[71][47]=1;ram[71][48]=1;ram[71][49]=1;ram[71][50]=1;ram[71][51]=1;ram[71][52]=1;ram[71][53]=1;ram[71][54]=0;ram[71][55]=1;ram[71][56]=1;ram[71][57]=1;ram[71][58]=1;ram[71][59]=0;ram[71][60]=0;ram[71][61]=1;ram[71][62]=1;ram[71][63]=1;ram[71][64]=0;ram[71][65]=0;ram[71][66]=0;ram[71][67]=0;ram[71][68]=0;ram[71][69]=1;ram[71][70]=0;ram[71][71]=1;ram[71][72]=1;ram[71][73]=1;ram[71][74]=1;ram[71][75]=0;ram[71][76]=1;ram[71][77]=1;ram[71][78]=0;ram[71][79]=1;ram[71][80]=0;ram[71][81]=1;ram[71][82]=0;ram[71][83]=1;ram[71][84]=0;ram[71][85]=0;ram[71][86]=0;ram[71][87]=0;ram[71][88]=1;ram[71][89]=1;ram[71][90]=1;ram[71][91]=0;ram[71][92]=0;ram[71][93]=1;ram[71][94]=0;ram[71][95]=1;ram[71][96]=1;ram[71][97]=1;ram[71][98]=0;ram[71][99]=0;ram[71][100]=0;ram[71][101]=1;ram[71][102]=0;ram[71][103]=1;ram[71][104]=1;ram[71][105]=1;ram[71][106]=1;ram[71][107]=1;ram[71][108]=1;ram[71][109]=1;ram[71][110]=1;ram[71][111]=0;ram[71][112]=1;ram[71][113]=1;ram[71][114]=0;ram[71][115]=0;ram[71][116]=0;ram[71][117]=1;ram[71][118]=0;ram[71][119]=1;ram[71][120]=1;ram[71][121]=0;ram[71][122]=0;ram[71][123]=1;ram[71][124]=1;ram[71][125]=0;ram[71][126]=1;ram[71][127]=1;ram[71][128]=1;ram[71][129]=1;ram[71][130]=1;ram[71][131]=1;ram[71][132]=0;ram[71][133]=1;ram[71][134]=1;ram[71][135]=1;ram[71][136]=0;
        ram[72][0]=1;ram[72][1]=0;ram[72][2]=0;ram[72][3]=1;ram[72][4]=1;ram[72][5]=1;ram[72][6]=1;ram[72][7]=1;ram[72][8]=0;ram[72][9]=0;ram[72][10]=1;ram[72][11]=0;ram[72][12]=1;ram[72][13]=0;ram[72][14]=0;ram[72][15]=1;ram[72][16]=1;ram[72][17]=1;ram[72][18]=1;ram[72][19]=1;ram[72][20]=1;ram[72][21]=0;ram[72][22]=0;ram[72][23]=1;ram[72][24]=1;ram[72][25]=1;ram[72][26]=1;ram[72][27]=0;ram[72][28]=1;ram[72][29]=1;ram[72][30]=1;ram[72][31]=1;ram[72][32]=1;ram[72][33]=1;ram[72][34]=1;ram[72][35]=1;ram[72][36]=1;ram[72][37]=1;ram[72][38]=1;ram[72][39]=1;ram[72][40]=1;ram[72][41]=0;ram[72][42]=0;ram[72][43]=1;ram[72][44]=0;ram[72][45]=1;ram[72][46]=1;ram[72][47]=1;ram[72][48]=1;ram[72][49]=0;ram[72][50]=0;ram[72][51]=0;ram[72][52]=1;ram[72][53]=1;ram[72][54]=1;ram[72][55]=1;ram[72][56]=1;ram[72][57]=1;ram[72][58]=1;ram[72][59]=0;ram[72][60]=1;ram[72][61]=0;ram[72][62]=1;ram[72][63]=1;ram[72][64]=1;ram[72][65]=1;ram[72][66]=1;ram[72][67]=1;ram[72][68]=1;ram[72][69]=0;ram[72][70]=1;ram[72][71]=0;ram[72][72]=1;ram[72][73]=1;ram[72][74]=0;ram[72][75]=1;ram[72][76]=1;ram[72][77]=0;ram[72][78]=1;ram[72][79]=0;ram[72][80]=0;ram[72][81]=1;ram[72][82]=0;ram[72][83]=0;ram[72][84]=1;ram[72][85]=1;ram[72][86]=1;ram[72][87]=1;ram[72][88]=1;ram[72][89]=1;ram[72][90]=0;ram[72][91]=0;ram[72][92]=0;ram[72][93]=1;ram[72][94]=1;ram[72][95]=1;ram[72][96]=0;ram[72][97]=1;ram[72][98]=1;ram[72][99]=1;ram[72][100]=0;ram[72][101]=1;ram[72][102]=1;ram[72][103]=1;ram[72][104]=1;ram[72][105]=0;ram[72][106]=1;ram[72][107]=1;ram[72][108]=1;ram[72][109]=1;ram[72][110]=1;ram[72][111]=0;ram[72][112]=0;ram[72][113]=1;ram[72][114]=1;ram[72][115]=1;ram[72][116]=0;ram[72][117]=1;ram[72][118]=0;ram[72][119]=1;ram[72][120]=0;ram[72][121]=0;ram[72][122]=0;ram[72][123]=1;ram[72][124]=1;ram[72][125]=1;ram[72][126]=1;ram[72][127]=0;ram[72][128]=0;ram[72][129]=1;ram[72][130]=0;ram[72][131]=1;ram[72][132]=1;ram[72][133]=0;ram[72][134]=1;ram[72][135]=0;ram[72][136]=1;
        ram[73][0]=1;ram[73][1]=1;ram[73][2]=0;ram[73][3]=0;ram[73][4]=1;ram[73][5]=0;ram[73][6]=0;ram[73][7]=1;ram[73][8]=0;ram[73][9]=0;ram[73][10]=1;ram[73][11]=1;ram[73][12]=1;ram[73][13]=1;ram[73][14]=0;ram[73][15]=1;ram[73][16]=0;ram[73][17]=1;ram[73][18]=0;ram[73][19]=1;ram[73][20]=1;ram[73][21]=1;ram[73][22]=1;ram[73][23]=1;ram[73][24]=1;ram[73][25]=1;ram[73][26]=1;ram[73][27]=1;ram[73][28]=0;ram[73][29]=1;ram[73][30]=1;ram[73][31]=1;ram[73][32]=1;ram[73][33]=1;ram[73][34]=0;ram[73][35]=1;ram[73][36]=0;ram[73][37]=1;ram[73][38]=1;ram[73][39]=1;ram[73][40]=0;ram[73][41]=1;ram[73][42]=1;ram[73][43]=0;ram[73][44]=1;ram[73][45]=1;ram[73][46]=0;ram[73][47]=1;ram[73][48]=1;ram[73][49]=0;ram[73][50]=0;ram[73][51]=1;ram[73][52]=0;ram[73][53]=1;ram[73][54]=0;ram[73][55]=0;ram[73][56]=1;ram[73][57]=0;ram[73][58]=1;ram[73][59]=1;ram[73][60]=1;ram[73][61]=1;ram[73][62]=1;ram[73][63]=1;ram[73][64]=1;ram[73][65]=0;ram[73][66]=1;ram[73][67]=0;ram[73][68]=0;ram[73][69]=1;ram[73][70]=0;ram[73][71]=1;ram[73][72]=1;ram[73][73]=0;ram[73][74]=1;ram[73][75]=1;ram[73][76]=1;ram[73][77]=0;ram[73][78]=1;ram[73][79]=0;ram[73][80]=0;ram[73][81]=0;ram[73][82]=1;ram[73][83]=0;ram[73][84]=1;ram[73][85]=0;ram[73][86]=1;ram[73][87]=1;ram[73][88]=1;ram[73][89]=1;ram[73][90]=0;ram[73][91]=1;ram[73][92]=0;ram[73][93]=1;ram[73][94]=1;ram[73][95]=1;ram[73][96]=0;ram[73][97]=1;ram[73][98]=1;ram[73][99]=1;ram[73][100]=1;ram[73][101]=1;ram[73][102]=1;ram[73][103]=1;ram[73][104]=1;ram[73][105]=1;ram[73][106]=1;ram[73][107]=0;ram[73][108]=0;ram[73][109]=0;ram[73][110]=0;ram[73][111]=0;ram[73][112]=0;ram[73][113]=1;ram[73][114]=1;ram[73][115]=0;ram[73][116]=1;ram[73][117]=1;ram[73][118]=0;ram[73][119]=1;ram[73][120]=0;ram[73][121]=0;ram[73][122]=1;ram[73][123]=0;ram[73][124]=1;ram[73][125]=0;ram[73][126]=0;ram[73][127]=1;ram[73][128]=0;ram[73][129]=0;ram[73][130]=1;ram[73][131]=1;ram[73][132]=0;ram[73][133]=1;ram[73][134]=1;ram[73][135]=1;ram[73][136]=1;
        ram[74][0]=1;ram[74][1]=0;ram[74][2]=1;ram[74][3]=0;ram[74][4]=1;ram[74][5]=1;ram[74][6]=0;ram[74][7]=0;ram[74][8]=1;ram[74][9]=1;ram[74][10]=1;ram[74][11]=1;ram[74][12]=1;ram[74][13]=1;ram[74][14]=0;ram[74][15]=1;ram[74][16]=1;ram[74][17]=0;ram[74][18]=0;ram[74][19]=1;ram[74][20]=0;ram[74][21]=1;ram[74][22]=1;ram[74][23]=1;ram[74][24]=0;ram[74][25]=1;ram[74][26]=1;ram[74][27]=1;ram[74][28]=1;ram[74][29]=0;ram[74][30]=1;ram[74][31]=1;ram[74][32]=0;ram[74][33]=0;ram[74][34]=1;ram[74][35]=0;ram[74][36]=1;ram[74][37]=0;ram[74][38]=1;ram[74][39]=1;ram[74][40]=1;ram[74][41]=0;ram[74][42]=0;ram[74][43]=1;ram[74][44]=0;ram[74][45]=0;ram[74][46]=0;ram[74][47]=0;ram[74][48]=1;ram[74][49]=1;ram[74][50]=0;ram[74][51]=0;ram[74][52]=1;ram[74][53]=0;ram[74][54]=0;ram[74][55]=0;ram[74][56]=1;ram[74][57]=1;ram[74][58]=1;ram[74][59]=1;ram[74][60]=1;ram[74][61]=1;ram[74][62]=1;ram[74][63]=1;ram[74][64]=1;ram[74][65]=1;ram[74][66]=0;ram[74][67]=1;ram[74][68]=1;ram[74][69]=1;ram[74][70]=0;ram[74][71]=0;ram[74][72]=1;ram[74][73]=0;ram[74][74]=0;ram[74][75]=1;ram[74][76]=0;ram[74][77]=1;ram[74][78]=1;ram[74][79]=1;ram[74][80]=1;ram[74][81]=1;ram[74][82]=1;ram[74][83]=1;ram[74][84]=1;ram[74][85]=1;ram[74][86]=1;ram[74][87]=0;ram[74][88]=1;ram[74][89]=0;ram[74][90]=1;ram[74][91]=1;ram[74][92]=1;ram[74][93]=1;ram[74][94]=1;ram[74][95]=0;ram[74][96]=1;ram[74][97]=1;ram[74][98]=0;ram[74][99]=1;ram[74][100]=0;ram[74][101]=0;ram[74][102]=0;ram[74][103]=1;ram[74][104]=0;ram[74][105]=1;ram[74][106]=1;ram[74][107]=1;ram[74][108]=0;ram[74][109]=0;ram[74][110]=1;ram[74][111]=1;ram[74][112]=0;ram[74][113]=1;ram[74][114]=0;ram[74][115]=0;ram[74][116]=1;ram[74][117]=0;ram[74][118]=1;ram[74][119]=1;ram[74][120]=1;ram[74][121]=1;ram[74][122]=0;ram[74][123]=1;ram[74][124]=0;ram[74][125]=1;ram[74][126]=1;ram[74][127]=1;ram[74][128]=1;ram[74][129]=1;ram[74][130]=1;ram[74][131]=1;ram[74][132]=0;ram[74][133]=1;ram[74][134]=1;ram[74][135]=0;ram[74][136]=1;
        ram[75][0]=1;ram[75][1]=1;ram[75][2]=1;ram[75][3]=1;ram[75][4]=0;ram[75][5]=1;ram[75][6]=0;ram[75][7]=0;ram[75][8]=1;ram[75][9]=1;ram[75][10]=1;ram[75][11]=1;ram[75][12]=1;ram[75][13]=1;ram[75][14]=1;ram[75][15]=0;ram[75][16]=1;ram[75][17]=1;ram[75][18]=1;ram[75][19]=0;ram[75][20]=1;ram[75][21]=0;ram[75][22]=1;ram[75][23]=0;ram[75][24]=1;ram[75][25]=1;ram[75][26]=1;ram[75][27]=0;ram[75][28]=0;ram[75][29]=1;ram[75][30]=0;ram[75][31]=1;ram[75][32]=1;ram[75][33]=0;ram[75][34]=1;ram[75][35]=1;ram[75][36]=1;ram[75][37]=1;ram[75][38]=0;ram[75][39]=1;ram[75][40]=0;ram[75][41]=1;ram[75][42]=1;ram[75][43]=1;ram[75][44]=0;ram[75][45]=1;ram[75][46]=1;ram[75][47]=0;ram[75][48]=1;ram[75][49]=1;ram[75][50]=1;ram[75][51]=0;ram[75][52]=1;ram[75][53]=1;ram[75][54]=1;ram[75][55]=1;ram[75][56]=0;ram[75][57]=1;ram[75][58]=0;ram[75][59]=1;ram[75][60]=1;ram[75][61]=0;ram[75][62]=1;ram[75][63]=0;ram[75][64]=0;ram[75][65]=1;ram[75][66]=1;ram[75][67]=1;ram[75][68]=1;ram[75][69]=0;ram[75][70]=1;ram[75][71]=1;ram[75][72]=1;ram[75][73]=1;ram[75][74]=1;ram[75][75]=1;ram[75][76]=1;ram[75][77]=0;ram[75][78]=0;ram[75][79]=1;ram[75][80]=1;ram[75][81]=0;ram[75][82]=1;ram[75][83]=1;ram[75][84]=1;ram[75][85]=1;ram[75][86]=1;ram[75][87]=0;ram[75][88]=1;ram[75][89]=1;ram[75][90]=1;ram[75][91]=0;ram[75][92]=0;ram[75][93]=0;ram[75][94]=1;ram[75][95]=0;ram[75][96]=1;ram[75][97]=0;ram[75][98]=0;ram[75][99]=0;ram[75][100]=0;ram[75][101]=1;ram[75][102]=1;ram[75][103]=1;ram[75][104]=0;ram[75][105]=0;ram[75][106]=0;ram[75][107]=0;ram[75][108]=0;ram[75][109]=1;ram[75][110]=1;ram[75][111]=1;ram[75][112]=1;ram[75][113]=1;ram[75][114]=1;ram[75][115]=1;ram[75][116]=1;ram[75][117]=0;ram[75][118]=1;ram[75][119]=1;ram[75][120]=1;ram[75][121]=1;ram[75][122]=0;ram[75][123]=0;ram[75][124]=0;ram[75][125]=1;ram[75][126]=1;ram[75][127]=0;ram[75][128]=0;ram[75][129]=1;ram[75][130]=1;ram[75][131]=0;ram[75][132]=1;ram[75][133]=0;ram[75][134]=1;ram[75][135]=1;ram[75][136]=1;
        ram[76][0]=0;ram[76][1]=1;ram[76][2]=0;ram[76][3]=1;ram[76][4]=0;ram[76][5]=0;ram[76][6]=1;ram[76][7]=1;ram[76][8]=0;ram[76][9]=1;ram[76][10]=0;ram[76][11]=1;ram[76][12]=1;ram[76][13]=1;ram[76][14]=0;ram[76][15]=0;ram[76][16]=1;ram[76][17]=1;ram[76][18]=1;ram[76][19]=0;ram[76][20]=0;ram[76][21]=1;ram[76][22]=1;ram[76][23]=1;ram[76][24]=1;ram[76][25]=1;ram[76][26]=1;ram[76][27]=1;ram[76][28]=0;ram[76][29]=0;ram[76][30]=1;ram[76][31]=1;ram[76][32]=0;ram[76][33]=0;ram[76][34]=0;ram[76][35]=0;ram[76][36]=1;ram[76][37]=1;ram[76][38]=1;ram[76][39]=0;ram[76][40]=1;ram[76][41]=1;ram[76][42]=0;ram[76][43]=1;ram[76][44]=1;ram[76][45]=1;ram[76][46]=0;ram[76][47]=1;ram[76][48]=1;ram[76][49]=1;ram[76][50]=0;ram[76][51]=1;ram[76][52]=0;ram[76][53]=1;ram[76][54]=1;ram[76][55]=0;ram[76][56]=1;ram[76][57]=1;ram[76][58]=1;ram[76][59]=1;ram[76][60]=1;ram[76][61]=1;ram[76][62]=1;ram[76][63]=1;ram[76][64]=1;ram[76][65]=1;ram[76][66]=1;ram[76][67]=1;ram[76][68]=1;ram[76][69]=1;ram[76][70]=1;ram[76][71]=1;ram[76][72]=1;ram[76][73]=1;ram[76][74]=1;ram[76][75]=1;ram[76][76]=1;ram[76][77]=1;ram[76][78]=1;ram[76][79]=1;ram[76][80]=1;ram[76][81]=0;ram[76][82]=1;ram[76][83]=0;ram[76][84]=1;ram[76][85]=1;ram[76][86]=1;ram[76][87]=1;ram[76][88]=1;ram[76][89]=1;ram[76][90]=1;ram[76][91]=1;ram[76][92]=1;ram[76][93]=1;ram[76][94]=1;ram[76][95]=1;ram[76][96]=0;ram[76][97]=1;ram[76][98]=1;ram[76][99]=1;ram[76][100]=0;ram[76][101]=1;ram[76][102]=0;ram[76][103]=1;ram[76][104]=1;ram[76][105]=0;ram[76][106]=1;ram[76][107]=1;ram[76][108]=1;ram[76][109]=1;ram[76][110]=1;ram[76][111]=1;ram[76][112]=1;ram[76][113]=1;ram[76][114]=1;ram[76][115]=0;ram[76][116]=1;ram[76][117]=1;ram[76][118]=0;ram[76][119]=1;ram[76][120]=1;ram[76][121]=1;ram[76][122]=1;ram[76][123]=0;ram[76][124]=1;ram[76][125]=1;ram[76][126]=0;ram[76][127]=1;ram[76][128]=0;ram[76][129]=1;ram[76][130]=0;ram[76][131]=1;ram[76][132]=1;ram[76][133]=1;ram[76][134]=1;ram[76][135]=1;ram[76][136]=1;
        ram[77][0]=1;ram[77][1]=1;ram[77][2]=1;ram[77][3]=0;ram[77][4]=0;ram[77][5]=1;ram[77][6]=1;ram[77][7]=0;ram[77][8]=1;ram[77][9]=1;ram[77][10]=0;ram[77][11]=1;ram[77][12]=0;ram[77][13]=1;ram[77][14]=1;ram[77][15]=1;ram[77][16]=0;ram[77][17]=1;ram[77][18]=1;ram[77][19]=0;ram[77][20]=0;ram[77][21]=1;ram[77][22]=1;ram[77][23]=0;ram[77][24]=1;ram[77][25]=0;ram[77][26]=0;ram[77][27]=1;ram[77][28]=1;ram[77][29]=0;ram[77][30]=0;ram[77][31]=1;ram[77][32]=1;ram[77][33]=0;ram[77][34]=0;ram[77][35]=1;ram[77][36]=0;ram[77][37]=1;ram[77][38]=1;ram[77][39]=1;ram[77][40]=1;ram[77][41]=1;ram[77][42]=1;ram[77][43]=1;ram[77][44]=1;ram[77][45]=1;ram[77][46]=0;ram[77][47]=1;ram[77][48]=1;ram[77][49]=0;ram[77][50]=1;ram[77][51]=1;ram[77][52]=1;ram[77][53]=1;ram[77][54]=1;ram[77][55]=1;ram[77][56]=0;ram[77][57]=1;ram[77][58]=1;ram[77][59]=1;ram[77][60]=1;ram[77][61]=0;ram[77][62]=1;ram[77][63]=0;ram[77][64]=1;ram[77][65]=1;ram[77][66]=0;ram[77][67]=1;ram[77][68]=0;ram[77][69]=1;ram[77][70]=1;ram[77][71]=1;ram[77][72]=1;ram[77][73]=0;ram[77][74]=0;ram[77][75]=1;ram[77][76]=1;ram[77][77]=1;ram[77][78]=1;ram[77][79]=0;ram[77][80]=1;ram[77][81]=1;ram[77][82]=1;ram[77][83]=0;ram[77][84]=1;ram[77][85]=1;ram[77][86]=1;ram[77][87]=1;ram[77][88]=1;ram[77][89]=1;ram[77][90]=1;ram[77][91]=0;ram[77][92]=1;ram[77][93]=1;ram[77][94]=1;ram[77][95]=1;ram[77][96]=1;ram[77][97]=1;ram[77][98]=0;ram[77][99]=1;ram[77][100]=1;ram[77][101]=1;ram[77][102]=0;ram[77][103]=1;ram[77][104]=1;ram[77][105]=0;ram[77][106]=0;ram[77][107]=1;ram[77][108]=1;ram[77][109]=1;ram[77][110]=1;ram[77][111]=0;ram[77][112]=0;ram[77][113]=1;ram[77][114]=1;ram[77][115]=0;ram[77][116]=0;ram[77][117]=1;ram[77][118]=1;ram[77][119]=1;ram[77][120]=0;ram[77][121]=0;ram[77][122]=0;ram[77][123]=1;ram[77][124]=1;ram[77][125]=1;ram[77][126]=1;ram[77][127]=0;ram[77][128]=0;ram[77][129]=1;ram[77][130]=1;ram[77][131]=0;ram[77][132]=0;ram[77][133]=0;ram[77][134]=0;ram[77][135]=0;ram[77][136]=1;
        ram[78][0]=1;ram[78][1]=0;ram[78][2]=1;ram[78][3]=1;ram[78][4]=1;ram[78][5]=1;ram[78][6]=1;ram[78][7]=0;ram[78][8]=0;ram[78][9]=0;ram[78][10]=1;ram[78][11]=1;ram[78][12]=1;ram[78][13]=0;ram[78][14]=0;ram[78][15]=1;ram[78][16]=1;ram[78][17]=0;ram[78][18]=1;ram[78][19]=0;ram[78][20]=1;ram[78][21]=1;ram[78][22]=1;ram[78][23]=0;ram[78][24]=1;ram[78][25]=0;ram[78][26]=1;ram[78][27]=1;ram[78][28]=0;ram[78][29]=0;ram[78][30]=1;ram[78][31]=1;ram[78][32]=0;ram[78][33]=1;ram[78][34]=0;ram[78][35]=1;ram[78][36]=1;ram[78][37]=1;ram[78][38]=1;ram[78][39]=1;ram[78][40]=1;ram[78][41]=0;ram[78][42]=0;ram[78][43]=0;ram[78][44]=0;ram[78][45]=1;ram[78][46]=1;ram[78][47]=0;ram[78][48]=1;ram[78][49]=0;ram[78][50]=1;ram[78][51]=0;ram[78][52]=1;ram[78][53]=1;ram[78][54]=1;ram[78][55]=1;ram[78][56]=0;ram[78][57]=1;ram[78][58]=1;ram[78][59]=0;ram[78][60]=1;ram[78][61]=1;ram[78][62]=1;ram[78][63]=1;ram[78][64]=1;ram[78][65]=1;ram[78][66]=1;ram[78][67]=1;ram[78][68]=0;ram[78][69]=1;ram[78][70]=0;ram[78][71]=0;ram[78][72]=0;ram[78][73]=1;ram[78][74]=1;ram[78][75]=1;ram[78][76]=0;ram[78][77]=0;ram[78][78]=1;ram[78][79]=1;ram[78][80]=0;ram[78][81]=0;ram[78][82]=1;ram[78][83]=0;ram[78][84]=1;ram[78][85]=1;ram[78][86]=1;ram[78][87]=1;ram[78][88]=1;ram[78][89]=1;ram[78][90]=0;ram[78][91]=1;ram[78][92]=0;ram[78][93]=0;ram[78][94]=1;ram[78][95]=0;ram[78][96]=1;ram[78][97]=1;ram[78][98]=0;ram[78][99]=1;ram[78][100]=1;ram[78][101]=1;ram[78][102]=1;ram[78][103]=1;ram[78][104]=1;ram[78][105]=1;ram[78][106]=1;ram[78][107]=1;ram[78][108]=0;ram[78][109]=0;ram[78][110]=0;ram[78][111]=1;ram[78][112]=1;ram[78][113]=0;ram[78][114]=1;ram[78][115]=1;ram[78][116]=1;ram[78][117]=1;ram[78][118]=1;ram[78][119]=1;ram[78][120]=1;ram[78][121]=0;ram[78][122]=1;ram[78][123]=1;ram[78][124]=0;ram[78][125]=0;ram[78][126]=0;ram[78][127]=1;ram[78][128]=0;ram[78][129]=1;ram[78][130]=1;ram[78][131]=0;ram[78][132]=1;ram[78][133]=1;ram[78][134]=1;ram[78][135]=1;ram[78][136]=1;
        ram[79][0]=1;ram[79][1]=1;ram[79][2]=1;ram[79][3]=1;ram[79][4]=0;ram[79][5]=1;ram[79][6]=1;ram[79][7]=1;ram[79][8]=0;ram[79][9]=1;ram[79][10]=0;ram[79][11]=0;ram[79][12]=0;ram[79][13]=1;ram[79][14]=1;ram[79][15]=0;ram[79][16]=1;ram[79][17]=1;ram[79][18]=1;ram[79][19]=0;ram[79][20]=0;ram[79][21]=1;ram[79][22]=0;ram[79][23]=1;ram[79][24]=1;ram[79][25]=1;ram[79][26]=0;ram[79][27]=1;ram[79][28]=1;ram[79][29]=1;ram[79][30]=1;ram[79][31]=0;ram[79][32]=0;ram[79][33]=1;ram[79][34]=0;ram[79][35]=1;ram[79][36]=1;ram[79][37]=0;ram[79][38]=1;ram[79][39]=1;ram[79][40]=0;ram[79][41]=0;ram[79][42]=1;ram[79][43]=0;ram[79][44]=1;ram[79][45]=1;ram[79][46]=1;ram[79][47]=0;ram[79][48]=1;ram[79][49]=1;ram[79][50]=1;ram[79][51]=1;ram[79][52]=1;ram[79][53]=1;ram[79][54]=0;ram[79][55]=0;ram[79][56]=1;ram[79][57]=1;ram[79][58]=1;ram[79][59]=1;ram[79][60]=1;ram[79][61]=0;ram[79][62]=0;ram[79][63]=1;ram[79][64]=1;ram[79][65]=1;ram[79][66]=0;ram[79][67]=1;ram[79][68]=1;ram[79][69]=0;ram[79][70]=0;ram[79][71]=1;ram[79][72]=1;ram[79][73]=0;ram[79][74]=0;ram[79][75]=1;ram[79][76]=1;ram[79][77]=1;ram[79][78]=1;ram[79][79]=1;ram[79][80]=1;ram[79][81]=1;ram[79][82]=1;ram[79][83]=1;ram[79][84]=1;ram[79][85]=0;ram[79][86]=1;ram[79][87]=0;ram[79][88]=1;ram[79][89]=1;ram[79][90]=0;ram[79][91]=1;ram[79][92]=0;ram[79][93]=0;ram[79][94]=1;ram[79][95]=1;ram[79][96]=1;ram[79][97]=1;ram[79][98]=1;ram[79][99]=1;ram[79][100]=0;ram[79][101]=1;ram[79][102]=1;ram[79][103]=1;ram[79][104]=1;ram[79][105]=1;ram[79][106]=0;ram[79][107]=1;ram[79][108]=1;ram[79][109]=0;ram[79][110]=1;ram[79][111]=1;ram[79][112]=0;ram[79][113]=0;ram[79][114]=1;ram[79][115]=1;ram[79][116]=0;ram[79][117]=1;ram[79][118]=0;ram[79][119]=0;ram[79][120]=0;ram[79][121]=1;ram[79][122]=1;ram[79][123]=1;ram[79][124]=0;ram[79][125]=1;ram[79][126]=1;ram[79][127]=1;ram[79][128]=1;ram[79][129]=1;ram[79][130]=1;ram[79][131]=0;ram[79][132]=1;ram[79][133]=1;ram[79][134]=1;ram[79][135]=1;ram[79][136]=0;
        ram[80][0]=0;ram[80][1]=1;ram[80][2]=1;ram[80][3]=1;ram[80][4]=0;ram[80][5]=0;ram[80][6]=1;ram[80][7]=0;ram[80][8]=1;ram[80][9]=1;ram[80][10]=0;ram[80][11]=0;ram[80][12]=0;ram[80][13]=0;ram[80][14]=0;ram[80][15]=1;ram[80][16]=1;ram[80][17]=1;ram[80][18]=1;ram[80][19]=1;ram[80][20]=1;ram[80][21]=1;ram[80][22]=1;ram[80][23]=1;ram[80][24]=1;ram[80][25]=0;ram[80][26]=1;ram[80][27]=1;ram[80][28]=1;ram[80][29]=1;ram[80][30]=1;ram[80][31]=0;ram[80][32]=1;ram[80][33]=1;ram[80][34]=1;ram[80][35]=1;ram[80][36]=1;ram[80][37]=1;ram[80][38]=0;ram[80][39]=0;ram[80][40]=1;ram[80][41]=0;ram[80][42]=1;ram[80][43]=1;ram[80][44]=1;ram[80][45]=0;ram[80][46]=0;ram[80][47]=0;ram[80][48]=0;ram[80][49]=1;ram[80][50]=1;ram[80][51]=1;ram[80][52]=1;ram[80][53]=1;ram[80][54]=0;ram[80][55]=1;ram[80][56]=0;ram[80][57]=1;ram[80][58]=0;ram[80][59]=1;ram[80][60]=1;ram[80][61]=1;ram[80][62]=1;ram[80][63]=0;ram[80][64]=0;ram[80][65]=0;ram[80][66]=1;ram[80][67]=0;ram[80][68]=1;ram[80][69]=1;ram[80][70]=1;ram[80][71]=1;ram[80][72]=0;ram[80][73]=1;ram[80][74]=1;ram[80][75]=1;ram[80][76]=1;ram[80][77]=1;ram[80][78]=1;ram[80][79]=0;ram[80][80]=1;ram[80][81]=0;ram[80][82]=1;ram[80][83]=1;ram[80][84]=1;ram[80][85]=1;ram[80][86]=0;ram[80][87]=1;ram[80][88]=1;ram[80][89]=1;ram[80][90]=1;ram[80][91]=1;ram[80][92]=1;ram[80][93]=0;ram[80][94]=0;ram[80][95]=0;ram[80][96]=0;ram[80][97]=0;ram[80][98]=0;ram[80][99]=0;ram[80][100]=1;ram[80][101]=0;ram[80][102]=0;ram[80][103]=0;ram[80][104]=0;ram[80][105]=0;ram[80][106]=1;ram[80][107]=1;ram[80][108]=1;ram[80][109]=1;ram[80][110]=1;ram[80][111]=0;ram[80][112]=0;ram[80][113]=0;ram[80][114]=0;ram[80][115]=0;ram[80][116]=1;ram[80][117]=1;ram[80][118]=0;ram[80][119]=1;ram[80][120]=1;ram[80][121]=0;ram[80][122]=1;ram[80][123]=0;ram[80][124]=1;ram[80][125]=1;ram[80][126]=1;ram[80][127]=1;ram[80][128]=0;ram[80][129]=1;ram[80][130]=1;ram[80][131]=0;ram[80][132]=0;ram[80][133]=0;ram[80][134]=0;ram[80][135]=1;ram[80][136]=1;
        ram[81][0]=0;ram[81][1]=1;ram[81][2]=1;ram[81][3]=1;ram[81][4]=1;ram[81][5]=0;ram[81][6]=0;ram[81][7]=1;ram[81][8]=0;ram[81][9]=1;ram[81][10]=1;ram[81][11]=1;ram[81][12]=1;ram[81][13]=0;ram[81][14]=0;ram[81][15]=0;ram[81][16]=1;ram[81][17]=0;ram[81][18]=1;ram[81][19]=0;ram[81][20]=1;ram[81][21]=0;ram[81][22]=0;ram[81][23]=1;ram[81][24]=1;ram[81][25]=1;ram[81][26]=0;ram[81][27]=0;ram[81][28]=1;ram[81][29]=1;ram[81][30]=0;ram[81][31]=1;ram[81][32]=1;ram[81][33]=1;ram[81][34]=0;ram[81][35]=1;ram[81][36]=1;ram[81][37]=0;ram[81][38]=1;ram[81][39]=1;ram[81][40]=0;ram[81][41]=1;ram[81][42]=0;ram[81][43]=1;ram[81][44]=0;ram[81][45]=0;ram[81][46]=0;ram[81][47]=1;ram[81][48]=0;ram[81][49]=0;ram[81][50]=1;ram[81][51]=0;ram[81][52]=1;ram[81][53]=0;ram[81][54]=1;ram[81][55]=1;ram[81][56]=1;ram[81][57]=1;ram[81][58]=1;ram[81][59]=0;ram[81][60]=1;ram[81][61]=1;ram[81][62]=1;ram[81][63]=1;ram[81][64]=1;ram[81][65]=0;ram[81][66]=1;ram[81][67]=1;ram[81][68]=1;ram[81][69]=0;ram[81][70]=1;ram[81][71]=0;ram[81][72]=1;ram[81][73]=1;ram[81][74]=1;ram[81][75]=0;ram[81][76]=1;ram[81][77]=1;ram[81][78]=1;ram[81][79]=0;ram[81][80]=1;ram[81][81]=1;ram[81][82]=1;ram[81][83]=0;ram[81][84]=1;ram[81][85]=0;ram[81][86]=1;ram[81][87]=1;ram[81][88]=1;ram[81][89]=1;ram[81][90]=0;ram[81][91]=0;ram[81][92]=1;ram[81][93]=1;ram[81][94]=0;ram[81][95]=0;ram[81][96]=1;ram[81][97]=1;ram[81][98]=1;ram[81][99]=0;ram[81][100]=0;ram[81][101]=1;ram[81][102]=1;ram[81][103]=0;ram[81][104]=1;ram[81][105]=1;ram[81][106]=0;ram[81][107]=0;ram[81][108]=1;ram[81][109]=1;ram[81][110]=0;ram[81][111]=1;ram[81][112]=1;ram[81][113]=1;ram[81][114]=1;ram[81][115]=0;ram[81][116]=1;ram[81][117]=1;ram[81][118]=0;ram[81][119]=1;ram[81][120]=1;ram[81][121]=1;ram[81][122]=1;ram[81][123]=1;ram[81][124]=1;ram[81][125]=1;ram[81][126]=1;ram[81][127]=1;ram[81][128]=0;ram[81][129]=0;ram[81][130]=0;ram[81][131]=1;ram[81][132]=1;ram[81][133]=1;ram[81][134]=0;ram[81][135]=1;ram[81][136]=1;
        ram[82][0]=0;ram[82][1]=1;ram[82][2]=1;ram[82][3]=1;ram[82][4]=0;ram[82][5]=1;ram[82][6]=1;ram[82][7]=0;ram[82][8]=1;ram[82][9]=1;ram[82][10]=1;ram[82][11]=1;ram[82][12]=1;ram[82][13]=1;ram[82][14]=0;ram[82][15]=0;ram[82][16]=0;ram[82][17]=0;ram[82][18]=0;ram[82][19]=1;ram[82][20]=0;ram[82][21]=0;ram[82][22]=0;ram[82][23]=0;ram[82][24]=1;ram[82][25]=1;ram[82][26]=1;ram[82][27]=0;ram[82][28]=1;ram[82][29]=1;ram[82][30]=0;ram[82][31]=0;ram[82][32]=0;ram[82][33]=0;ram[82][34]=1;ram[82][35]=1;ram[82][36]=0;ram[82][37]=1;ram[82][38]=1;ram[82][39]=1;ram[82][40]=1;ram[82][41]=1;ram[82][42]=1;ram[82][43]=0;ram[82][44]=0;ram[82][45]=1;ram[82][46]=1;ram[82][47]=0;ram[82][48]=1;ram[82][49]=1;ram[82][50]=1;ram[82][51]=1;ram[82][52]=1;ram[82][53]=1;ram[82][54]=1;ram[82][55]=1;ram[82][56]=1;ram[82][57]=1;ram[82][58]=1;ram[82][59]=1;ram[82][60]=0;ram[82][61]=1;ram[82][62]=1;ram[82][63]=1;ram[82][64]=0;ram[82][65]=1;ram[82][66]=0;ram[82][67]=0;ram[82][68]=1;ram[82][69]=1;ram[82][70]=0;ram[82][71]=1;ram[82][72]=1;ram[82][73]=1;ram[82][74]=1;ram[82][75]=1;ram[82][76]=0;ram[82][77]=1;ram[82][78]=1;ram[82][79]=1;ram[82][80]=1;ram[82][81]=1;ram[82][82]=0;ram[82][83]=0;ram[82][84]=0;ram[82][85]=0;ram[82][86]=1;ram[82][87]=1;ram[82][88]=0;ram[82][89]=1;ram[82][90]=1;ram[82][91]=0;ram[82][92]=1;ram[82][93]=1;ram[82][94]=1;ram[82][95]=0;ram[82][96]=1;ram[82][97]=1;ram[82][98]=1;ram[82][99]=0;ram[82][100]=1;ram[82][101]=0;ram[82][102]=0;ram[82][103]=0;ram[82][104]=1;ram[82][105]=1;ram[82][106]=1;ram[82][107]=1;ram[82][108]=1;ram[82][109]=1;ram[82][110]=0;ram[82][111]=1;ram[82][112]=0;ram[82][113]=0;ram[82][114]=1;ram[82][115]=1;ram[82][116]=1;ram[82][117]=1;ram[82][118]=1;ram[82][119]=1;ram[82][120]=0;ram[82][121]=0;ram[82][122]=0;ram[82][123]=1;ram[82][124]=0;ram[82][125]=1;ram[82][126]=0;ram[82][127]=0;ram[82][128]=1;ram[82][129]=1;ram[82][130]=1;ram[82][131]=0;ram[82][132]=1;ram[82][133]=1;ram[82][134]=1;ram[82][135]=0;ram[82][136]=1;
        ram[83][0]=0;ram[83][1]=1;ram[83][2]=1;ram[83][3]=1;ram[83][4]=0;ram[83][5]=0;ram[83][6]=1;ram[83][7]=0;ram[83][8]=1;ram[83][9]=1;ram[83][10]=1;ram[83][11]=0;ram[83][12]=0;ram[83][13]=0;ram[83][14]=1;ram[83][15]=0;ram[83][16]=1;ram[83][17]=1;ram[83][18]=0;ram[83][19]=0;ram[83][20]=0;ram[83][21]=1;ram[83][22]=0;ram[83][23]=1;ram[83][24]=0;ram[83][25]=0;ram[83][26]=1;ram[83][27]=0;ram[83][28]=1;ram[83][29]=0;ram[83][30]=0;ram[83][31]=1;ram[83][32]=0;ram[83][33]=0;ram[83][34]=1;ram[83][35]=0;ram[83][36]=0;ram[83][37]=0;ram[83][38]=0;ram[83][39]=1;ram[83][40]=1;ram[83][41]=1;ram[83][42]=0;ram[83][43]=0;ram[83][44]=0;ram[83][45]=1;ram[83][46]=1;ram[83][47]=1;ram[83][48]=1;ram[83][49]=1;ram[83][50]=1;ram[83][51]=0;ram[83][52]=1;ram[83][53]=0;ram[83][54]=1;ram[83][55]=1;ram[83][56]=0;ram[83][57]=1;ram[83][58]=1;ram[83][59]=1;ram[83][60]=1;ram[83][61]=1;ram[83][62]=1;ram[83][63]=0;ram[83][64]=0;ram[83][65]=1;ram[83][66]=1;ram[83][67]=1;ram[83][68]=1;ram[83][69]=0;ram[83][70]=0;ram[83][71]=1;ram[83][72]=1;ram[83][73]=1;ram[83][74]=1;ram[83][75]=1;ram[83][76]=1;ram[83][77]=1;ram[83][78]=1;ram[83][79]=1;ram[83][80]=0;ram[83][81]=1;ram[83][82]=0;ram[83][83]=0;ram[83][84]=1;ram[83][85]=1;ram[83][86]=1;ram[83][87]=1;ram[83][88]=0;ram[83][89]=0;ram[83][90]=1;ram[83][91]=1;ram[83][92]=1;ram[83][93]=1;ram[83][94]=1;ram[83][95]=1;ram[83][96]=0;ram[83][97]=0;ram[83][98]=1;ram[83][99]=1;ram[83][100]=1;ram[83][101]=0;ram[83][102]=1;ram[83][103]=1;ram[83][104]=0;ram[83][105]=1;ram[83][106]=0;ram[83][107]=1;ram[83][108]=1;ram[83][109]=0;ram[83][110]=1;ram[83][111]=1;ram[83][112]=1;ram[83][113]=0;ram[83][114]=1;ram[83][115]=0;ram[83][116]=0;ram[83][117]=0;ram[83][118]=0;ram[83][119]=0;ram[83][120]=0;ram[83][121]=0;ram[83][122]=1;ram[83][123]=1;ram[83][124]=1;ram[83][125]=1;ram[83][126]=0;ram[83][127]=1;ram[83][128]=0;ram[83][129]=0;ram[83][130]=0;ram[83][131]=1;ram[83][132]=1;ram[83][133]=0;ram[83][134]=0;ram[83][135]=1;ram[83][136]=1;
        ram[84][0]=1;ram[84][1]=1;ram[84][2]=1;ram[84][3]=1;ram[84][4]=0;ram[84][5]=0;ram[84][6]=1;ram[84][7]=1;ram[84][8]=0;ram[84][9]=1;ram[84][10]=0;ram[84][11]=0;ram[84][12]=1;ram[84][13]=0;ram[84][14]=1;ram[84][15]=0;ram[84][16]=1;ram[84][17]=1;ram[84][18]=0;ram[84][19]=1;ram[84][20]=1;ram[84][21]=0;ram[84][22]=0;ram[84][23]=0;ram[84][24]=1;ram[84][25]=0;ram[84][26]=1;ram[84][27]=1;ram[84][28]=0;ram[84][29]=1;ram[84][30]=0;ram[84][31]=0;ram[84][32]=0;ram[84][33]=0;ram[84][34]=1;ram[84][35]=1;ram[84][36]=1;ram[84][37]=1;ram[84][38]=0;ram[84][39]=1;ram[84][40]=0;ram[84][41]=1;ram[84][42]=0;ram[84][43]=1;ram[84][44]=0;ram[84][45]=1;ram[84][46]=0;ram[84][47]=0;ram[84][48]=1;ram[84][49]=0;ram[84][50]=1;ram[84][51]=1;ram[84][52]=1;ram[84][53]=1;ram[84][54]=0;ram[84][55]=0;ram[84][56]=1;ram[84][57]=0;ram[84][58]=1;ram[84][59]=1;ram[84][60]=1;ram[84][61]=1;ram[84][62]=0;ram[84][63]=1;ram[84][64]=1;ram[84][65]=1;ram[84][66]=1;ram[84][67]=1;ram[84][68]=1;ram[84][69]=1;ram[84][70]=1;ram[84][71]=0;ram[84][72]=0;ram[84][73]=1;ram[84][74]=1;ram[84][75]=0;ram[84][76]=0;ram[84][77]=1;ram[84][78]=1;ram[84][79]=1;ram[84][80]=1;ram[84][81]=1;ram[84][82]=1;ram[84][83]=0;ram[84][84]=0;ram[84][85]=1;ram[84][86]=1;ram[84][87]=1;ram[84][88]=0;ram[84][89]=1;ram[84][90]=1;ram[84][91]=1;ram[84][92]=1;ram[84][93]=1;ram[84][94]=0;ram[84][95]=0;ram[84][96]=1;ram[84][97]=1;ram[84][98]=1;ram[84][99]=0;ram[84][100]=1;ram[84][101]=0;ram[84][102]=0;ram[84][103]=1;ram[84][104]=1;ram[84][105]=1;ram[84][106]=1;ram[84][107]=1;ram[84][108]=1;ram[84][109]=0;ram[84][110]=1;ram[84][111]=1;ram[84][112]=0;ram[84][113]=0;ram[84][114]=1;ram[84][115]=1;ram[84][116]=1;ram[84][117]=1;ram[84][118]=0;ram[84][119]=0;ram[84][120]=0;ram[84][121]=1;ram[84][122]=0;ram[84][123]=1;ram[84][124]=1;ram[84][125]=0;ram[84][126]=1;ram[84][127]=0;ram[84][128]=0;ram[84][129]=1;ram[84][130]=0;ram[84][131]=0;ram[84][132]=0;ram[84][133]=0;ram[84][134]=1;ram[84][135]=1;ram[84][136]=0;
        ram[85][0]=1;ram[85][1]=0;ram[85][2]=1;ram[85][3]=1;ram[85][4]=0;ram[85][5]=1;ram[85][6]=0;ram[85][7]=0;ram[85][8]=1;ram[85][9]=1;ram[85][10]=0;ram[85][11]=1;ram[85][12]=0;ram[85][13]=0;ram[85][14]=0;ram[85][15]=0;ram[85][16]=0;ram[85][17]=1;ram[85][18]=1;ram[85][19]=0;ram[85][20]=1;ram[85][21]=1;ram[85][22]=1;ram[85][23]=0;ram[85][24]=1;ram[85][25]=0;ram[85][26]=1;ram[85][27]=0;ram[85][28]=1;ram[85][29]=0;ram[85][30]=1;ram[85][31]=1;ram[85][32]=1;ram[85][33]=1;ram[85][34]=0;ram[85][35]=1;ram[85][36]=1;ram[85][37]=0;ram[85][38]=1;ram[85][39]=1;ram[85][40]=1;ram[85][41]=0;ram[85][42]=0;ram[85][43]=1;ram[85][44]=0;ram[85][45]=0;ram[85][46]=0;ram[85][47]=1;ram[85][48]=1;ram[85][49]=0;ram[85][50]=1;ram[85][51]=1;ram[85][52]=0;ram[85][53]=1;ram[85][54]=0;ram[85][55]=1;ram[85][56]=0;ram[85][57]=0;ram[85][58]=1;ram[85][59]=1;ram[85][60]=1;ram[85][61]=1;ram[85][62]=0;ram[85][63]=0;ram[85][64]=0;ram[85][65]=0;ram[85][66]=0;ram[85][67]=1;ram[85][68]=1;ram[85][69]=1;ram[85][70]=1;ram[85][71]=0;ram[85][72]=0;ram[85][73]=1;ram[85][74]=1;ram[85][75]=1;ram[85][76]=0;ram[85][77]=1;ram[85][78]=0;ram[85][79]=1;ram[85][80]=1;ram[85][81]=0;ram[85][82]=1;ram[85][83]=0;ram[85][84]=1;ram[85][85]=1;ram[85][86]=1;ram[85][87]=0;ram[85][88]=1;ram[85][89]=0;ram[85][90]=1;ram[85][91]=1;ram[85][92]=1;ram[85][93]=0;ram[85][94]=1;ram[85][95]=1;ram[85][96]=1;ram[85][97]=1;ram[85][98]=0;ram[85][99]=1;ram[85][100]=1;ram[85][101]=0;ram[85][102]=1;ram[85][103]=1;ram[85][104]=1;ram[85][105]=1;ram[85][106]=1;ram[85][107]=1;ram[85][108]=0;ram[85][109]=1;ram[85][110]=0;ram[85][111]=1;ram[85][112]=1;ram[85][113]=0;ram[85][114]=1;ram[85][115]=0;ram[85][116]=1;ram[85][117]=1;ram[85][118]=0;ram[85][119]=1;ram[85][120]=1;ram[85][121]=0;ram[85][122]=1;ram[85][123]=1;ram[85][124]=1;ram[85][125]=1;ram[85][126]=0;ram[85][127]=1;ram[85][128]=0;ram[85][129]=0;ram[85][130]=1;ram[85][131]=0;ram[85][132]=0;ram[85][133]=1;ram[85][134]=0;ram[85][135]=1;ram[85][136]=1;
        ram[86][0]=0;ram[86][1]=1;ram[86][2]=0;ram[86][3]=1;ram[86][4]=0;ram[86][5]=0;ram[86][6]=1;ram[86][7]=1;ram[86][8]=1;ram[86][9]=1;ram[86][10]=0;ram[86][11]=1;ram[86][12]=1;ram[86][13]=0;ram[86][14]=0;ram[86][15]=1;ram[86][16]=1;ram[86][17]=1;ram[86][18]=0;ram[86][19]=0;ram[86][20]=0;ram[86][21]=1;ram[86][22]=1;ram[86][23]=1;ram[86][24]=1;ram[86][25]=0;ram[86][26]=0;ram[86][27]=0;ram[86][28]=1;ram[86][29]=1;ram[86][30]=1;ram[86][31]=1;ram[86][32]=0;ram[86][33]=1;ram[86][34]=0;ram[86][35]=0;ram[86][36]=1;ram[86][37]=1;ram[86][38]=1;ram[86][39]=1;ram[86][40]=1;ram[86][41]=1;ram[86][42]=0;ram[86][43]=1;ram[86][44]=0;ram[86][45]=0;ram[86][46]=0;ram[86][47]=1;ram[86][48]=1;ram[86][49]=1;ram[86][50]=0;ram[86][51]=0;ram[86][52]=1;ram[86][53]=0;ram[86][54]=1;ram[86][55]=1;ram[86][56]=0;ram[86][57]=0;ram[86][58]=0;ram[86][59]=1;ram[86][60]=1;ram[86][61]=1;ram[86][62]=0;ram[86][63]=1;ram[86][64]=1;ram[86][65]=1;ram[86][66]=1;ram[86][67]=1;ram[86][68]=0;ram[86][69]=0;ram[86][70]=1;ram[86][71]=1;ram[86][72]=0;ram[86][73]=0;ram[86][74]=0;ram[86][75]=0;ram[86][76]=1;ram[86][77]=1;ram[86][78]=0;ram[86][79]=1;ram[86][80]=1;ram[86][81]=1;ram[86][82]=1;ram[86][83]=1;ram[86][84]=1;ram[86][85]=1;ram[86][86]=1;ram[86][87]=0;ram[86][88]=0;ram[86][89]=1;ram[86][90]=0;ram[86][91]=1;ram[86][92]=0;ram[86][93]=1;ram[86][94]=0;ram[86][95]=1;ram[86][96]=0;ram[86][97]=1;ram[86][98]=1;ram[86][99]=1;ram[86][100]=1;ram[86][101]=0;ram[86][102]=1;ram[86][103]=1;ram[86][104]=1;ram[86][105]=0;ram[86][106]=0;ram[86][107]=1;ram[86][108]=1;ram[86][109]=1;ram[86][110]=1;ram[86][111]=0;ram[86][112]=1;ram[86][113]=1;ram[86][114]=1;ram[86][115]=1;ram[86][116]=1;ram[86][117]=1;ram[86][118]=0;ram[86][119]=0;ram[86][120]=1;ram[86][121]=0;ram[86][122]=1;ram[86][123]=1;ram[86][124]=0;ram[86][125]=1;ram[86][126]=0;ram[86][127]=1;ram[86][128]=1;ram[86][129]=0;ram[86][130]=1;ram[86][131]=1;ram[86][132]=1;ram[86][133]=1;ram[86][134]=0;ram[86][135]=1;ram[86][136]=1;
        ram[87][0]=1;ram[87][1]=0;ram[87][2]=0;ram[87][3]=1;ram[87][4]=1;ram[87][5]=0;ram[87][6]=0;ram[87][7]=0;ram[87][8]=1;ram[87][9]=0;ram[87][10]=1;ram[87][11]=0;ram[87][12]=0;ram[87][13]=0;ram[87][14]=1;ram[87][15]=0;ram[87][16]=0;ram[87][17]=0;ram[87][18]=0;ram[87][19]=1;ram[87][20]=1;ram[87][21]=1;ram[87][22]=1;ram[87][23]=1;ram[87][24]=0;ram[87][25]=1;ram[87][26]=1;ram[87][27]=1;ram[87][28]=0;ram[87][29]=1;ram[87][30]=0;ram[87][31]=0;ram[87][32]=0;ram[87][33]=1;ram[87][34]=0;ram[87][35]=0;ram[87][36]=0;ram[87][37]=1;ram[87][38]=0;ram[87][39]=0;ram[87][40]=1;ram[87][41]=1;ram[87][42]=1;ram[87][43]=0;ram[87][44]=1;ram[87][45]=1;ram[87][46]=1;ram[87][47]=1;ram[87][48]=0;ram[87][49]=0;ram[87][50]=0;ram[87][51]=1;ram[87][52]=1;ram[87][53]=1;ram[87][54]=1;ram[87][55]=1;ram[87][56]=1;ram[87][57]=1;ram[87][58]=0;ram[87][59]=1;ram[87][60]=1;ram[87][61]=1;ram[87][62]=1;ram[87][63]=1;ram[87][64]=1;ram[87][65]=0;ram[87][66]=1;ram[87][67]=1;ram[87][68]=1;ram[87][69]=0;ram[87][70]=1;ram[87][71]=1;ram[87][72]=1;ram[87][73]=1;ram[87][74]=1;ram[87][75]=0;ram[87][76]=1;ram[87][77]=0;ram[87][78]=0;ram[87][79]=0;ram[87][80]=1;ram[87][81]=0;ram[87][82]=0;ram[87][83]=1;ram[87][84]=1;ram[87][85]=1;ram[87][86]=0;ram[87][87]=1;ram[87][88]=0;ram[87][89]=1;ram[87][90]=1;ram[87][91]=0;ram[87][92]=1;ram[87][93]=1;ram[87][94]=1;ram[87][95]=0;ram[87][96]=0;ram[87][97]=1;ram[87][98]=1;ram[87][99]=1;ram[87][100]=1;ram[87][101]=0;ram[87][102]=0;ram[87][103]=0;ram[87][104]=1;ram[87][105]=1;ram[87][106]=0;ram[87][107]=0;ram[87][108]=0;ram[87][109]=1;ram[87][110]=1;ram[87][111]=1;ram[87][112]=0;ram[87][113]=1;ram[87][114]=0;ram[87][115]=0;ram[87][116]=0;ram[87][117]=1;ram[87][118]=1;ram[87][119]=0;ram[87][120]=1;ram[87][121]=1;ram[87][122]=0;ram[87][123]=1;ram[87][124]=0;ram[87][125]=1;ram[87][126]=1;ram[87][127]=0;ram[87][128]=0;ram[87][129]=1;ram[87][130]=0;ram[87][131]=1;ram[87][132]=1;ram[87][133]=1;ram[87][134]=1;ram[87][135]=0;ram[87][136]=0;
        ram[88][0]=1;ram[88][1]=1;ram[88][2]=1;ram[88][3]=1;ram[88][4]=1;ram[88][5]=1;ram[88][6]=1;ram[88][7]=0;ram[88][8]=0;ram[88][9]=0;ram[88][10]=1;ram[88][11]=1;ram[88][12]=1;ram[88][13]=1;ram[88][14]=1;ram[88][15]=0;ram[88][16]=1;ram[88][17]=0;ram[88][18]=0;ram[88][19]=0;ram[88][20]=0;ram[88][21]=1;ram[88][22]=1;ram[88][23]=0;ram[88][24]=1;ram[88][25]=1;ram[88][26]=0;ram[88][27]=0;ram[88][28]=1;ram[88][29]=0;ram[88][30]=1;ram[88][31]=1;ram[88][32]=1;ram[88][33]=1;ram[88][34]=0;ram[88][35]=0;ram[88][36]=1;ram[88][37]=1;ram[88][38]=0;ram[88][39]=0;ram[88][40]=1;ram[88][41]=0;ram[88][42]=0;ram[88][43]=0;ram[88][44]=1;ram[88][45]=1;ram[88][46]=0;ram[88][47]=1;ram[88][48]=1;ram[88][49]=1;ram[88][50]=1;ram[88][51]=1;ram[88][52]=0;ram[88][53]=1;ram[88][54]=1;ram[88][55]=0;ram[88][56]=0;ram[88][57]=1;ram[88][58]=1;ram[88][59]=0;ram[88][60]=0;ram[88][61]=1;ram[88][62]=1;ram[88][63]=1;ram[88][64]=0;ram[88][65]=0;ram[88][66]=1;ram[88][67]=0;ram[88][68]=1;ram[88][69]=1;ram[88][70]=0;ram[88][71]=1;ram[88][72]=0;ram[88][73]=1;ram[88][74]=0;ram[88][75]=0;ram[88][76]=1;ram[88][77]=0;ram[88][78]=0;ram[88][79]=1;ram[88][80]=1;ram[88][81]=0;ram[88][82]=0;ram[88][83]=0;ram[88][84]=1;ram[88][85]=1;ram[88][86]=1;ram[88][87]=0;ram[88][88]=0;ram[88][89]=1;ram[88][90]=0;ram[88][91]=1;ram[88][92]=1;ram[88][93]=1;ram[88][94]=1;ram[88][95]=1;ram[88][96]=0;ram[88][97]=0;ram[88][98]=0;ram[88][99]=1;ram[88][100]=0;ram[88][101]=0;ram[88][102]=1;ram[88][103]=0;ram[88][104]=1;ram[88][105]=1;ram[88][106]=1;ram[88][107]=1;ram[88][108]=1;ram[88][109]=1;ram[88][110]=1;ram[88][111]=1;ram[88][112]=1;ram[88][113]=1;ram[88][114]=0;ram[88][115]=0;ram[88][116]=1;ram[88][117]=0;ram[88][118]=0;ram[88][119]=1;ram[88][120]=0;ram[88][121]=1;ram[88][122]=0;ram[88][123]=1;ram[88][124]=1;ram[88][125]=0;ram[88][126]=1;ram[88][127]=1;ram[88][128]=0;ram[88][129]=1;ram[88][130]=0;ram[88][131]=1;ram[88][132]=0;ram[88][133]=1;ram[88][134]=1;ram[88][135]=0;ram[88][136]=1;
        ram[89][0]=1;ram[89][1]=1;ram[89][2]=1;ram[89][3]=0;ram[89][4]=1;ram[89][5]=1;ram[89][6]=0;ram[89][7]=0;ram[89][8]=1;ram[89][9]=1;ram[89][10]=1;ram[89][11]=0;ram[89][12]=1;ram[89][13]=1;ram[89][14]=1;ram[89][15]=1;ram[89][16]=0;ram[89][17]=1;ram[89][18]=1;ram[89][19]=1;ram[89][20]=1;ram[89][21]=1;ram[89][22]=1;ram[89][23]=0;ram[89][24]=0;ram[89][25]=0;ram[89][26]=1;ram[89][27]=1;ram[89][28]=0;ram[89][29]=0;ram[89][30]=1;ram[89][31]=0;ram[89][32]=1;ram[89][33]=1;ram[89][34]=1;ram[89][35]=1;ram[89][36]=1;ram[89][37]=0;ram[89][38]=0;ram[89][39]=1;ram[89][40]=1;ram[89][41]=1;ram[89][42]=1;ram[89][43]=0;ram[89][44]=0;ram[89][45]=1;ram[89][46]=0;ram[89][47]=1;ram[89][48]=1;ram[89][49]=1;ram[89][50]=1;ram[89][51]=1;ram[89][52]=0;ram[89][53]=1;ram[89][54]=1;ram[89][55]=0;ram[89][56]=0;ram[89][57]=0;ram[89][58]=0;ram[89][59]=0;ram[89][60]=1;ram[89][61]=1;ram[89][62]=1;ram[89][63]=0;ram[89][64]=0;ram[89][65]=1;ram[89][66]=0;ram[89][67]=1;ram[89][68]=1;ram[89][69]=1;ram[89][70]=1;ram[89][71]=0;ram[89][72]=0;ram[89][73]=1;ram[89][74]=0;ram[89][75]=1;ram[89][76]=0;ram[89][77]=0;ram[89][78]=1;ram[89][79]=0;ram[89][80]=1;ram[89][81]=1;ram[89][82]=1;ram[89][83]=1;ram[89][84]=1;ram[89][85]=1;ram[89][86]=0;ram[89][87]=0;ram[89][88]=1;ram[89][89]=1;ram[89][90]=0;ram[89][91]=1;ram[89][92]=1;ram[89][93]=1;ram[89][94]=0;ram[89][95]=1;ram[89][96]=0;ram[89][97]=1;ram[89][98]=0;ram[89][99]=0;ram[89][100]=1;ram[89][101]=1;ram[89][102]=1;ram[89][103]=1;ram[89][104]=1;ram[89][105]=0;ram[89][106]=0;ram[89][107]=0;ram[89][108]=0;ram[89][109]=1;ram[89][110]=0;ram[89][111]=1;ram[89][112]=1;ram[89][113]=1;ram[89][114]=1;ram[89][115]=1;ram[89][116]=1;ram[89][117]=1;ram[89][118]=1;ram[89][119]=0;ram[89][120]=0;ram[89][121]=1;ram[89][122]=0;ram[89][123]=1;ram[89][124]=1;ram[89][125]=1;ram[89][126]=1;ram[89][127]=1;ram[89][128]=0;ram[89][129]=1;ram[89][130]=0;ram[89][131]=1;ram[89][132]=1;ram[89][133]=1;ram[89][134]=1;ram[89][135]=0;ram[89][136]=0;
        ram[90][0]=1;ram[90][1]=1;ram[90][2]=1;ram[90][3]=0;ram[90][4]=1;ram[90][5]=0;ram[90][6]=0;ram[90][7]=0;ram[90][8]=1;ram[90][9]=0;ram[90][10]=1;ram[90][11]=1;ram[90][12]=1;ram[90][13]=1;ram[90][14]=0;ram[90][15]=1;ram[90][16]=0;ram[90][17]=1;ram[90][18]=0;ram[90][19]=1;ram[90][20]=1;ram[90][21]=0;ram[90][22]=1;ram[90][23]=1;ram[90][24]=0;ram[90][25]=1;ram[90][26]=1;ram[90][27]=0;ram[90][28]=0;ram[90][29]=1;ram[90][30]=0;ram[90][31]=1;ram[90][32]=1;ram[90][33]=1;ram[90][34]=1;ram[90][35]=1;ram[90][36]=1;ram[90][37]=1;ram[90][38]=0;ram[90][39]=1;ram[90][40]=1;ram[90][41]=0;ram[90][42]=0;ram[90][43]=1;ram[90][44]=1;ram[90][45]=1;ram[90][46]=0;ram[90][47]=0;ram[90][48]=1;ram[90][49]=1;ram[90][50]=1;ram[90][51]=1;ram[90][52]=0;ram[90][53]=1;ram[90][54]=0;ram[90][55]=0;ram[90][56]=0;ram[90][57]=0;ram[90][58]=1;ram[90][59]=1;ram[90][60]=0;ram[90][61]=1;ram[90][62]=0;ram[90][63]=1;ram[90][64]=1;ram[90][65]=1;ram[90][66]=1;ram[90][67]=1;ram[90][68]=1;ram[90][69]=0;ram[90][70]=1;ram[90][71]=0;ram[90][72]=1;ram[90][73]=1;ram[90][74]=1;ram[90][75]=1;ram[90][76]=1;ram[90][77]=0;ram[90][78]=0;ram[90][79]=1;ram[90][80]=0;ram[90][81]=1;ram[90][82]=1;ram[90][83]=1;ram[90][84]=1;ram[90][85]=1;ram[90][86]=1;ram[90][87]=1;ram[90][88]=0;ram[90][89]=1;ram[90][90]=0;ram[90][91]=1;ram[90][92]=0;ram[90][93]=1;ram[90][94]=1;ram[90][95]=1;ram[90][96]=0;ram[90][97]=0;ram[90][98]=0;ram[90][99]=0;ram[90][100]=1;ram[90][101]=1;ram[90][102]=1;ram[90][103]=0;ram[90][104]=1;ram[90][105]=1;ram[90][106]=1;ram[90][107]=0;ram[90][108]=1;ram[90][109]=1;ram[90][110]=1;ram[90][111]=1;ram[90][112]=0;ram[90][113]=1;ram[90][114]=1;ram[90][115]=0;ram[90][116]=1;ram[90][117]=1;ram[90][118]=1;ram[90][119]=0;ram[90][120]=0;ram[90][121]=1;ram[90][122]=1;ram[90][123]=1;ram[90][124]=1;ram[90][125]=1;ram[90][126]=1;ram[90][127]=1;ram[90][128]=1;ram[90][129]=1;ram[90][130]=1;ram[90][131]=1;ram[90][132]=1;ram[90][133]=1;ram[90][134]=1;ram[90][135]=1;ram[90][136]=1;
        ram[91][0]=1;ram[91][1]=1;ram[91][2]=0;ram[91][3]=0;ram[91][4]=0;ram[91][5]=0;ram[91][6]=0;ram[91][7]=1;ram[91][8]=1;ram[91][9]=0;ram[91][10]=0;ram[91][11]=1;ram[91][12]=0;ram[91][13]=1;ram[91][14]=0;ram[91][15]=0;ram[91][16]=1;ram[91][17]=1;ram[91][18]=1;ram[91][19]=0;ram[91][20]=1;ram[91][21]=0;ram[91][22]=0;ram[91][23]=0;ram[91][24]=1;ram[91][25]=0;ram[91][26]=0;ram[91][27]=0;ram[91][28]=1;ram[91][29]=0;ram[91][30]=0;ram[91][31]=0;ram[91][32]=0;ram[91][33]=1;ram[91][34]=0;ram[91][35]=1;ram[91][36]=1;ram[91][37]=0;ram[91][38]=1;ram[91][39]=0;ram[91][40]=0;ram[91][41]=1;ram[91][42]=0;ram[91][43]=1;ram[91][44]=1;ram[91][45]=0;ram[91][46]=1;ram[91][47]=1;ram[91][48]=1;ram[91][49]=1;ram[91][50]=0;ram[91][51]=1;ram[91][52]=0;ram[91][53]=1;ram[91][54]=0;ram[91][55]=0;ram[91][56]=1;ram[91][57]=0;ram[91][58]=0;ram[91][59]=1;ram[91][60]=0;ram[91][61]=1;ram[91][62]=1;ram[91][63]=1;ram[91][64]=1;ram[91][65]=0;ram[91][66]=1;ram[91][67]=1;ram[91][68]=0;ram[91][69]=0;ram[91][70]=1;ram[91][71]=0;ram[91][72]=1;ram[91][73]=0;ram[91][74]=1;ram[91][75]=0;ram[91][76]=1;ram[91][77]=1;ram[91][78]=0;ram[91][79]=1;ram[91][80]=1;ram[91][81]=1;ram[91][82]=0;ram[91][83]=1;ram[91][84]=0;ram[91][85]=0;ram[91][86]=1;ram[91][87]=1;ram[91][88]=1;ram[91][89]=1;ram[91][90]=1;ram[91][91]=0;ram[91][92]=0;ram[91][93]=1;ram[91][94]=0;ram[91][95]=1;ram[91][96]=0;ram[91][97]=0;ram[91][98]=1;ram[91][99]=0;ram[91][100]=1;ram[91][101]=1;ram[91][102]=0;ram[91][103]=0;ram[91][104]=1;ram[91][105]=0;ram[91][106]=0;ram[91][107]=0;ram[91][108]=0;ram[91][109]=1;ram[91][110]=0;ram[91][111]=1;ram[91][112]=1;ram[91][113]=1;ram[91][114]=0;ram[91][115]=0;ram[91][116]=1;ram[91][117]=0;ram[91][118]=1;ram[91][119]=1;ram[91][120]=0;ram[91][121]=1;ram[91][122]=1;ram[91][123]=1;ram[91][124]=1;ram[91][125]=1;ram[91][126]=1;ram[91][127]=1;ram[91][128]=1;ram[91][129]=0;ram[91][130]=1;ram[91][131]=1;ram[91][132]=1;ram[91][133]=1;ram[91][134]=0;ram[91][135]=1;ram[91][136]=0;
        ram[92][0]=1;ram[92][1]=1;ram[92][2]=1;ram[92][3]=0;ram[92][4]=0;ram[92][5]=0;ram[92][6]=1;ram[92][7]=1;ram[92][8]=1;ram[92][9]=0;ram[92][10]=1;ram[92][11]=0;ram[92][12]=0;ram[92][13]=1;ram[92][14]=0;ram[92][15]=1;ram[92][16]=1;ram[92][17]=0;ram[92][18]=0;ram[92][19]=1;ram[92][20]=0;ram[92][21]=0;ram[92][22]=1;ram[92][23]=0;ram[92][24]=0;ram[92][25]=1;ram[92][26]=1;ram[92][27]=1;ram[92][28]=1;ram[92][29]=0;ram[92][30]=1;ram[92][31]=0;ram[92][32]=1;ram[92][33]=1;ram[92][34]=1;ram[92][35]=0;ram[92][36]=1;ram[92][37]=0;ram[92][38]=1;ram[92][39]=1;ram[92][40]=1;ram[92][41]=1;ram[92][42]=1;ram[92][43]=1;ram[92][44]=1;ram[92][45]=1;ram[92][46]=1;ram[92][47]=0;ram[92][48]=1;ram[92][49]=1;ram[92][50]=1;ram[92][51]=0;ram[92][52]=0;ram[92][53]=1;ram[92][54]=0;ram[92][55]=1;ram[92][56]=1;ram[92][57]=0;ram[92][58]=0;ram[92][59]=1;ram[92][60]=1;ram[92][61]=1;ram[92][62]=1;ram[92][63]=0;ram[92][64]=0;ram[92][65]=1;ram[92][66]=0;ram[92][67]=1;ram[92][68]=0;ram[92][69]=0;ram[92][70]=1;ram[92][71]=1;ram[92][72]=0;ram[92][73]=1;ram[92][74]=1;ram[92][75]=1;ram[92][76]=1;ram[92][77]=1;ram[92][78]=1;ram[92][79]=1;ram[92][80]=0;ram[92][81]=1;ram[92][82]=1;ram[92][83]=1;ram[92][84]=1;ram[92][85]=1;ram[92][86]=1;ram[92][87]=1;ram[92][88]=0;ram[92][89]=1;ram[92][90]=0;ram[92][91]=0;ram[92][92]=1;ram[92][93]=1;ram[92][94]=1;ram[92][95]=0;ram[92][96]=0;ram[92][97]=1;ram[92][98]=1;ram[92][99]=1;ram[92][100]=1;ram[92][101]=1;ram[92][102]=1;ram[92][103]=1;ram[92][104]=0;ram[92][105]=1;ram[92][106]=0;ram[92][107]=0;ram[92][108]=1;ram[92][109]=0;ram[92][110]=1;ram[92][111]=1;ram[92][112]=1;ram[92][113]=1;ram[92][114]=0;ram[92][115]=1;ram[92][116]=1;ram[92][117]=1;ram[92][118]=0;ram[92][119]=0;ram[92][120]=0;ram[92][121]=1;ram[92][122]=1;ram[92][123]=1;ram[92][124]=0;ram[92][125]=1;ram[92][126]=1;ram[92][127]=0;ram[92][128]=1;ram[92][129]=0;ram[92][130]=0;ram[92][131]=1;ram[92][132]=1;ram[92][133]=1;ram[92][134]=0;ram[92][135]=1;ram[92][136]=1;
        ram[93][0]=1;ram[93][1]=1;ram[93][2]=1;ram[93][3]=0;ram[93][4]=1;ram[93][5]=0;ram[93][6]=1;ram[93][7]=0;ram[93][8]=1;ram[93][9]=1;ram[93][10]=1;ram[93][11]=0;ram[93][12]=1;ram[93][13]=0;ram[93][14]=1;ram[93][15]=0;ram[93][16]=0;ram[93][17]=0;ram[93][18]=1;ram[93][19]=1;ram[93][20]=1;ram[93][21]=0;ram[93][22]=0;ram[93][23]=1;ram[93][24]=0;ram[93][25]=0;ram[93][26]=1;ram[93][27]=0;ram[93][28]=1;ram[93][29]=0;ram[93][30]=1;ram[93][31]=1;ram[93][32]=0;ram[93][33]=1;ram[93][34]=1;ram[93][35]=1;ram[93][36]=1;ram[93][37]=1;ram[93][38]=1;ram[93][39]=1;ram[93][40]=1;ram[93][41]=0;ram[93][42]=0;ram[93][43]=1;ram[93][44]=1;ram[93][45]=1;ram[93][46]=1;ram[93][47]=1;ram[93][48]=0;ram[93][49]=1;ram[93][50]=0;ram[93][51]=1;ram[93][52]=0;ram[93][53]=0;ram[93][54]=1;ram[93][55]=1;ram[93][56]=0;ram[93][57]=1;ram[93][58]=0;ram[93][59]=1;ram[93][60]=1;ram[93][61]=0;ram[93][62]=1;ram[93][63]=1;ram[93][64]=1;ram[93][65]=0;ram[93][66]=1;ram[93][67]=0;ram[93][68]=1;ram[93][69]=1;ram[93][70]=0;ram[93][71]=0;ram[93][72]=1;ram[93][73]=0;ram[93][74]=1;ram[93][75]=1;ram[93][76]=1;ram[93][77]=1;ram[93][78]=1;ram[93][79]=1;ram[93][80]=0;ram[93][81]=1;ram[93][82]=0;ram[93][83]=1;ram[93][84]=0;ram[93][85]=1;ram[93][86]=1;ram[93][87]=0;ram[93][88]=0;ram[93][89]=0;ram[93][90]=0;ram[93][91]=0;ram[93][92]=1;ram[93][93]=0;ram[93][94]=0;ram[93][95]=0;ram[93][96]=1;ram[93][97]=1;ram[93][98]=1;ram[93][99]=1;ram[93][100]=1;ram[93][101]=1;ram[93][102]=1;ram[93][103]=1;ram[93][104]=1;ram[93][105]=0;ram[93][106]=1;ram[93][107]=1;ram[93][108]=0;ram[93][109]=1;ram[93][110]=0;ram[93][111]=1;ram[93][112]=0;ram[93][113]=1;ram[93][114]=1;ram[93][115]=1;ram[93][116]=1;ram[93][117]=0;ram[93][118]=1;ram[93][119]=1;ram[93][120]=0;ram[93][121]=1;ram[93][122]=1;ram[93][123]=0;ram[93][124]=1;ram[93][125]=0;ram[93][126]=1;ram[93][127]=1;ram[93][128]=1;ram[93][129]=1;ram[93][130]=1;ram[93][131]=0;ram[93][132]=0;ram[93][133]=0;ram[93][134]=1;ram[93][135]=0;ram[93][136]=1;
        ram[94][0]=1;ram[94][1]=1;ram[94][2]=1;ram[94][3]=0;ram[94][4]=1;ram[94][5]=0;ram[94][6]=1;ram[94][7]=0;ram[94][8]=1;ram[94][9]=1;ram[94][10]=0;ram[94][11]=0;ram[94][12]=1;ram[94][13]=1;ram[94][14]=0;ram[94][15]=1;ram[94][16]=1;ram[94][17]=1;ram[94][18]=1;ram[94][19]=1;ram[94][20]=0;ram[94][21]=1;ram[94][22]=1;ram[94][23]=1;ram[94][24]=1;ram[94][25]=0;ram[94][26]=0;ram[94][27]=1;ram[94][28]=1;ram[94][29]=1;ram[94][30]=1;ram[94][31]=1;ram[94][32]=1;ram[94][33]=1;ram[94][34]=0;ram[94][35]=0;ram[94][36]=0;ram[94][37]=1;ram[94][38]=0;ram[94][39]=0;ram[94][40]=0;ram[94][41]=1;ram[94][42]=0;ram[94][43]=1;ram[94][44]=0;ram[94][45]=1;ram[94][46]=1;ram[94][47]=1;ram[94][48]=0;ram[94][49]=0;ram[94][50]=1;ram[94][51]=1;ram[94][52]=1;ram[94][53]=1;ram[94][54]=1;ram[94][55]=1;ram[94][56]=0;ram[94][57]=1;ram[94][58]=1;ram[94][59]=1;ram[94][60]=1;ram[94][61]=0;ram[94][62]=0;ram[94][63]=1;ram[94][64]=1;ram[94][65]=1;ram[94][66]=0;ram[94][67]=1;ram[94][68]=0;ram[94][69]=0;ram[94][70]=1;ram[94][71]=0;ram[94][72]=1;ram[94][73]=0;ram[94][74]=1;ram[94][75]=1;ram[94][76]=1;ram[94][77]=0;ram[94][78]=1;ram[94][79]=0;ram[94][80]=0;ram[94][81]=1;ram[94][82]=0;ram[94][83]=1;ram[94][84]=1;ram[94][85]=1;ram[94][86]=1;ram[94][87]=1;ram[94][88]=0;ram[94][89]=1;ram[94][90]=1;ram[94][91]=1;ram[94][92]=1;ram[94][93]=0;ram[94][94]=0;ram[94][95]=1;ram[94][96]=1;ram[94][97]=1;ram[94][98]=1;ram[94][99]=0;ram[94][100]=1;ram[94][101]=1;ram[94][102]=1;ram[94][103]=1;ram[94][104]=0;ram[94][105]=0;ram[94][106]=1;ram[94][107]=0;ram[94][108]=1;ram[94][109]=0;ram[94][110]=1;ram[94][111]=0;ram[94][112]=1;ram[94][113]=1;ram[94][114]=1;ram[94][115]=0;ram[94][116]=1;ram[94][117]=1;ram[94][118]=1;ram[94][119]=1;ram[94][120]=0;ram[94][121]=1;ram[94][122]=1;ram[94][123]=1;ram[94][124]=1;ram[94][125]=1;ram[94][126]=1;ram[94][127]=0;ram[94][128]=0;ram[94][129]=1;ram[94][130]=0;ram[94][131]=1;ram[94][132]=1;ram[94][133]=1;ram[94][134]=1;ram[94][135]=0;ram[94][136]=1;
        ram[95][0]=1;ram[95][1]=1;ram[95][2]=1;ram[95][3]=1;ram[95][4]=0;ram[95][5]=1;ram[95][6]=0;ram[95][7]=1;ram[95][8]=1;ram[95][9]=1;ram[95][10]=1;ram[95][11]=1;ram[95][12]=1;ram[95][13]=0;ram[95][14]=1;ram[95][15]=1;ram[95][16]=1;ram[95][17]=1;ram[95][18]=1;ram[95][19]=1;ram[95][20]=0;ram[95][21]=0;ram[95][22]=0;ram[95][23]=0;ram[95][24]=0;ram[95][25]=1;ram[95][26]=0;ram[95][27]=1;ram[95][28]=0;ram[95][29]=1;ram[95][30]=1;ram[95][31]=1;ram[95][32]=0;ram[95][33]=1;ram[95][34]=0;ram[95][35]=1;ram[95][36]=1;ram[95][37]=1;ram[95][38]=1;ram[95][39]=0;ram[95][40]=1;ram[95][41]=1;ram[95][42]=1;ram[95][43]=1;ram[95][44]=1;ram[95][45]=1;ram[95][46]=1;ram[95][47]=0;ram[95][48]=1;ram[95][49]=1;ram[95][50]=0;ram[95][51]=0;ram[95][52]=1;ram[95][53]=1;ram[95][54]=1;ram[95][55]=1;ram[95][56]=1;ram[95][57]=1;ram[95][58]=1;ram[95][59]=1;ram[95][60]=1;ram[95][61]=1;ram[95][62]=1;ram[95][63]=1;ram[95][64]=0;ram[95][65]=0;ram[95][66]=0;ram[95][67]=0;ram[95][68]=1;ram[95][69]=1;ram[95][70]=1;ram[95][71]=1;ram[95][72]=0;ram[95][73]=0;ram[95][74]=0;ram[95][75]=1;ram[95][76]=0;ram[95][77]=1;ram[95][78]=0;ram[95][79]=1;ram[95][80]=0;ram[95][81]=1;ram[95][82]=1;ram[95][83]=0;ram[95][84]=1;ram[95][85]=0;ram[95][86]=1;ram[95][87]=0;ram[95][88]=1;ram[95][89]=0;ram[95][90]=1;ram[95][91]=0;ram[95][92]=0;ram[95][93]=0;ram[95][94]=0;ram[95][95]=0;ram[95][96]=1;ram[95][97]=1;ram[95][98]=0;ram[95][99]=1;ram[95][100]=1;ram[95][101]=1;ram[95][102]=1;ram[95][103]=0;ram[95][104]=1;ram[95][105]=0;ram[95][106]=1;ram[95][107]=1;ram[95][108]=0;ram[95][109]=0;ram[95][110]=0;ram[95][111]=1;ram[95][112]=0;ram[95][113]=0;ram[95][114]=0;ram[95][115]=0;ram[95][116]=1;ram[95][117]=1;ram[95][118]=1;ram[95][119]=1;ram[95][120]=1;ram[95][121]=0;ram[95][122]=0;ram[95][123]=1;ram[95][124]=1;ram[95][125]=0;ram[95][126]=0;ram[95][127]=0;ram[95][128]=1;ram[95][129]=1;ram[95][130]=1;ram[95][131]=1;ram[95][132]=1;ram[95][133]=1;ram[95][134]=0;ram[95][135]=1;ram[95][136]=0;
        ram[96][0]=1;ram[96][1]=0;ram[96][2]=1;ram[96][3]=1;ram[96][4]=1;ram[96][5]=0;ram[96][6]=1;ram[96][7]=1;ram[96][8]=0;ram[96][9]=1;ram[96][10]=1;ram[96][11]=1;ram[96][12]=1;ram[96][13]=0;ram[96][14]=1;ram[96][15]=1;ram[96][16]=0;ram[96][17]=1;ram[96][18]=0;ram[96][19]=0;ram[96][20]=1;ram[96][21]=1;ram[96][22]=0;ram[96][23]=1;ram[96][24]=1;ram[96][25]=1;ram[96][26]=1;ram[96][27]=0;ram[96][28]=0;ram[96][29]=1;ram[96][30]=1;ram[96][31]=1;ram[96][32]=1;ram[96][33]=1;ram[96][34]=1;ram[96][35]=0;ram[96][36]=1;ram[96][37]=0;ram[96][38]=1;ram[96][39]=0;ram[96][40]=0;ram[96][41]=1;ram[96][42]=1;ram[96][43]=1;ram[96][44]=1;ram[96][45]=1;ram[96][46]=1;ram[96][47]=0;ram[96][48]=0;ram[96][49]=1;ram[96][50]=0;ram[96][51]=1;ram[96][52]=0;ram[96][53]=1;ram[96][54]=0;ram[96][55]=1;ram[96][56]=1;ram[96][57]=0;ram[96][58]=1;ram[96][59]=1;ram[96][60]=0;ram[96][61]=0;ram[96][62]=1;ram[96][63]=1;ram[96][64]=1;ram[96][65]=1;ram[96][66]=1;ram[96][67]=0;ram[96][68]=1;ram[96][69]=1;ram[96][70]=1;ram[96][71]=1;ram[96][72]=0;ram[96][73]=0;ram[96][74]=0;ram[96][75]=1;ram[96][76]=1;ram[96][77]=1;ram[96][78]=1;ram[96][79]=1;ram[96][80]=0;ram[96][81]=1;ram[96][82]=1;ram[96][83]=1;ram[96][84]=1;ram[96][85]=0;ram[96][86]=1;ram[96][87]=1;ram[96][88]=1;ram[96][89]=1;ram[96][90]=1;ram[96][91]=1;ram[96][92]=1;ram[96][93]=0;ram[96][94]=0;ram[96][95]=0;ram[96][96]=1;ram[96][97]=0;ram[96][98]=1;ram[96][99]=1;ram[96][100]=0;ram[96][101]=1;ram[96][102]=1;ram[96][103]=1;ram[96][104]=1;ram[96][105]=1;ram[96][106]=0;ram[96][107]=0;ram[96][108]=0;ram[96][109]=1;ram[96][110]=1;ram[96][111]=1;ram[96][112]=1;ram[96][113]=1;ram[96][114]=1;ram[96][115]=1;ram[96][116]=1;ram[96][117]=1;ram[96][118]=1;ram[96][119]=1;ram[96][120]=1;ram[96][121]=0;ram[96][122]=1;ram[96][123]=1;ram[96][124]=1;ram[96][125]=1;ram[96][126]=1;ram[96][127]=0;ram[96][128]=0;ram[96][129]=1;ram[96][130]=0;ram[96][131]=1;ram[96][132]=0;ram[96][133]=0;ram[96][134]=1;ram[96][135]=1;ram[96][136]=1;
        ram[97][0]=0;ram[97][1]=1;ram[97][2]=0;ram[97][3]=0;ram[97][4]=0;ram[97][5]=0;ram[97][6]=0;ram[97][7]=1;ram[97][8]=1;ram[97][9]=0;ram[97][10]=0;ram[97][11]=1;ram[97][12]=1;ram[97][13]=0;ram[97][14]=1;ram[97][15]=0;ram[97][16]=1;ram[97][17]=1;ram[97][18]=1;ram[97][19]=1;ram[97][20]=0;ram[97][21]=1;ram[97][22]=1;ram[97][23]=0;ram[97][24]=1;ram[97][25]=0;ram[97][26]=1;ram[97][27]=1;ram[97][28]=0;ram[97][29]=1;ram[97][30]=1;ram[97][31]=0;ram[97][32]=1;ram[97][33]=0;ram[97][34]=1;ram[97][35]=1;ram[97][36]=1;ram[97][37]=1;ram[97][38]=1;ram[97][39]=0;ram[97][40]=1;ram[97][41]=0;ram[97][42]=1;ram[97][43]=0;ram[97][44]=1;ram[97][45]=1;ram[97][46]=0;ram[97][47]=1;ram[97][48]=0;ram[97][49]=1;ram[97][50]=1;ram[97][51]=1;ram[97][52]=1;ram[97][53]=0;ram[97][54]=1;ram[97][55]=1;ram[97][56]=1;ram[97][57]=1;ram[97][58]=0;ram[97][59]=0;ram[97][60]=0;ram[97][61]=1;ram[97][62]=0;ram[97][63]=1;ram[97][64]=1;ram[97][65]=1;ram[97][66]=1;ram[97][67]=1;ram[97][68]=1;ram[97][69]=1;ram[97][70]=0;ram[97][71]=0;ram[97][72]=1;ram[97][73]=1;ram[97][74]=1;ram[97][75]=0;ram[97][76]=0;ram[97][77]=1;ram[97][78]=1;ram[97][79]=1;ram[97][80]=1;ram[97][81]=1;ram[97][82]=0;ram[97][83]=1;ram[97][84]=1;ram[97][85]=1;ram[97][86]=1;ram[97][87]=0;ram[97][88]=1;ram[97][89]=0;ram[97][90]=1;ram[97][91]=0;ram[97][92]=1;ram[97][93]=0;ram[97][94]=1;ram[97][95]=0;ram[97][96]=0;ram[97][97]=0;ram[97][98]=1;ram[97][99]=0;ram[97][100]=0;ram[97][101]=0;ram[97][102]=1;ram[97][103]=0;ram[97][104]=1;ram[97][105]=1;ram[97][106]=0;ram[97][107]=1;ram[97][108]=1;ram[97][109]=1;ram[97][110]=0;ram[97][111]=0;ram[97][112]=0;ram[97][113]=1;ram[97][114]=1;ram[97][115]=0;ram[97][116]=0;ram[97][117]=1;ram[97][118]=1;ram[97][119]=1;ram[97][120]=0;ram[97][121]=1;ram[97][122]=0;ram[97][123]=1;ram[97][124]=1;ram[97][125]=1;ram[97][126]=1;ram[97][127]=1;ram[97][128]=0;ram[97][129]=1;ram[97][130]=0;ram[97][131]=0;ram[97][132]=1;ram[97][133]=1;ram[97][134]=1;ram[97][135]=0;ram[97][136]=1;
        ram[98][0]=1;ram[98][1]=1;ram[98][2]=1;ram[98][3]=1;ram[98][4]=0;ram[98][5]=1;ram[98][6]=1;ram[98][7]=0;ram[98][8]=0;ram[98][9]=0;ram[98][10]=0;ram[98][11]=0;ram[98][12]=1;ram[98][13]=1;ram[98][14]=0;ram[98][15]=1;ram[98][16]=0;ram[98][17]=1;ram[98][18]=0;ram[98][19]=1;ram[98][20]=1;ram[98][21]=1;ram[98][22]=0;ram[98][23]=1;ram[98][24]=0;ram[98][25]=1;ram[98][26]=0;ram[98][27]=1;ram[98][28]=1;ram[98][29]=1;ram[98][30]=1;ram[98][31]=1;ram[98][32]=0;ram[98][33]=1;ram[98][34]=1;ram[98][35]=1;ram[98][36]=0;ram[98][37]=0;ram[98][38]=0;ram[98][39]=1;ram[98][40]=1;ram[98][41]=1;ram[98][42]=1;ram[98][43]=1;ram[98][44]=1;ram[98][45]=1;ram[98][46]=0;ram[98][47]=1;ram[98][48]=0;ram[98][49]=1;ram[98][50]=1;ram[98][51]=1;ram[98][52]=0;ram[98][53]=1;ram[98][54]=0;ram[98][55]=0;ram[98][56]=0;ram[98][57]=1;ram[98][58]=0;ram[98][59]=1;ram[98][60]=1;ram[98][61]=1;ram[98][62]=1;ram[98][63]=0;ram[98][64]=1;ram[98][65]=1;ram[98][66]=1;ram[98][67]=1;ram[98][68]=1;ram[98][69]=1;ram[98][70]=1;ram[98][71]=1;ram[98][72]=0;ram[98][73]=1;ram[98][74]=1;ram[98][75]=1;ram[98][76]=1;ram[98][77]=1;ram[98][78]=1;ram[98][79]=0;ram[98][80]=0;ram[98][81]=0;ram[98][82]=0;ram[98][83]=1;ram[98][84]=1;ram[98][85]=1;ram[98][86]=1;ram[98][87]=0;ram[98][88]=1;ram[98][89]=1;ram[98][90]=1;ram[98][91]=0;ram[98][92]=0;ram[98][93]=1;ram[98][94]=1;ram[98][95]=0;ram[98][96]=1;ram[98][97]=1;ram[98][98]=1;ram[98][99]=0;ram[98][100]=0;ram[98][101]=1;ram[98][102]=1;ram[98][103]=1;ram[98][104]=1;ram[98][105]=0;ram[98][106]=1;ram[98][107]=1;ram[98][108]=0;ram[98][109]=1;ram[98][110]=1;ram[98][111]=1;ram[98][112]=0;ram[98][113]=0;ram[98][114]=1;ram[98][115]=0;ram[98][116]=1;ram[98][117]=1;ram[98][118]=0;ram[98][119]=1;ram[98][120]=1;ram[98][121]=0;ram[98][122]=1;ram[98][123]=1;ram[98][124]=1;ram[98][125]=1;ram[98][126]=1;ram[98][127]=1;ram[98][128]=1;ram[98][129]=1;ram[98][130]=1;ram[98][131]=1;ram[98][132]=0;ram[98][133]=0;ram[98][134]=1;ram[98][135]=1;ram[98][136]=0;
        ram[99][0]=0;ram[99][1]=1;ram[99][2]=1;ram[99][3]=1;ram[99][4]=1;ram[99][5]=1;ram[99][6]=1;ram[99][7]=1;ram[99][8]=0;ram[99][9]=1;ram[99][10]=1;ram[99][11]=1;ram[99][12]=1;ram[99][13]=0;ram[99][14]=1;ram[99][15]=0;ram[99][16]=1;ram[99][17]=1;ram[99][18]=0;ram[99][19]=0;ram[99][20]=1;ram[99][21]=1;ram[99][22]=1;ram[99][23]=1;ram[99][24]=1;ram[99][25]=1;ram[99][26]=1;ram[99][27]=1;ram[99][28]=1;ram[99][29]=0;ram[99][30]=1;ram[99][31]=1;ram[99][32]=1;ram[99][33]=1;ram[99][34]=1;ram[99][35]=0;ram[99][36]=0;ram[99][37]=0;ram[99][38]=0;ram[99][39]=1;ram[99][40]=0;ram[99][41]=0;ram[99][42]=1;ram[99][43]=0;ram[99][44]=0;ram[99][45]=1;ram[99][46]=1;ram[99][47]=0;ram[99][48]=1;ram[99][49]=1;ram[99][50]=1;ram[99][51]=1;ram[99][52]=1;ram[99][53]=1;ram[99][54]=1;ram[99][55]=0;ram[99][56]=0;ram[99][57]=1;ram[99][58]=0;ram[99][59]=0;ram[99][60]=1;ram[99][61]=1;ram[99][62]=1;ram[99][63]=0;ram[99][64]=0;ram[99][65]=0;ram[99][66]=1;ram[99][67]=1;ram[99][68]=1;ram[99][69]=1;ram[99][70]=1;ram[99][71]=1;ram[99][72]=0;ram[99][73]=1;ram[99][74]=1;ram[99][75]=0;ram[99][76]=1;ram[99][77]=1;ram[99][78]=0;ram[99][79]=0;ram[99][80]=1;ram[99][81]=1;ram[99][82]=1;ram[99][83]=1;ram[99][84]=1;ram[99][85]=0;ram[99][86]=0;ram[99][87]=0;ram[99][88]=1;ram[99][89]=1;ram[99][90]=1;ram[99][91]=1;ram[99][92]=0;ram[99][93]=1;ram[99][94]=1;ram[99][95]=1;ram[99][96]=1;ram[99][97]=0;ram[99][98]=0;ram[99][99]=1;ram[99][100]=0;ram[99][101]=1;ram[99][102]=0;ram[99][103]=1;ram[99][104]=1;ram[99][105]=1;ram[99][106]=1;ram[99][107]=0;ram[99][108]=0;ram[99][109]=1;ram[99][110]=1;ram[99][111]=1;ram[99][112]=1;ram[99][113]=0;ram[99][114]=0;ram[99][115]=1;ram[99][116]=0;ram[99][117]=0;ram[99][118]=0;ram[99][119]=1;ram[99][120]=1;ram[99][121]=0;ram[99][122]=1;ram[99][123]=1;ram[99][124]=1;ram[99][125]=1;ram[99][126]=1;ram[99][127]=1;ram[99][128]=1;ram[99][129]=0;ram[99][130]=1;ram[99][131]=1;ram[99][132]=0;ram[99][133]=0;ram[99][134]=0;ram[99][135]=0;ram[99][136]=0;
        ram[100][0]=1;ram[100][1]=0;ram[100][2]=1;ram[100][3]=0;ram[100][4]=1;ram[100][5]=0;ram[100][6]=1;ram[100][7]=1;ram[100][8]=1;ram[100][9]=1;ram[100][10]=1;ram[100][11]=1;ram[100][12]=1;ram[100][13]=0;ram[100][14]=0;ram[100][15]=0;ram[100][16]=1;ram[100][17]=1;ram[100][18]=0;ram[100][19]=1;ram[100][20]=1;ram[100][21]=1;ram[100][22]=0;ram[100][23]=0;ram[100][24]=0;ram[100][25]=1;ram[100][26]=0;ram[100][27]=1;ram[100][28]=1;ram[100][29]=0;ram[100][30]=1;ram[100][31]=0;ram[100][32]=0;ram[100][33]=1;ram[100][34]=0;ram[100][35]=1;ram[100][36]=0;ram[100][37]=1;ram[100][38]=0;ram[100][39]=1;ram[100][40]=1;ram[100][41]=1;ram[100][42]=0;ram[100][43]=1;ram[100][44]=1;ram[100][45]=0;ram[100][46]=0;ram[100][47]=1;ram[100][48]=1;ram[100][49]=1;ram[100][50]=0;ram[100][51]=1;ram[100][52]=1;ram[100][53]=1;ram[100][54]=1;ram[100][55]=0;ram[100][56]=0;ram[100][57]=1;ram[100][58]=0;ram[100][59]=0;ram[100][60]=0;ram[100][61]=0;ram[100][62]=1;ram[100][63]=0;ram[100][64]=0;ram[100][65]=1;ram[100][66]=1;ram[100][67]=1;ram[100][68]=0;ram[100][69]=1;ram[100][70]=0;ram[100][71]=0;ram[100][72]=1;ram[100][73]=0;ram[100][74]=1;ram[100][75]=0;ram[100][76]=0;ram[100][77]=0;ram[100][78]=0;ram[100][79]=1;ram[100][80]=0;ram[100][81]=1;ram[100][82]=1;ram[100][83]=1;ram[100][84]=0;ram[100][85]=1;ram[100][86]=0;ram[100][87]=1;ram[100][88]=0;ram[100][89]=1;ram[100][90]=1;ram[100][91]=0;ram[100][92]=1;ram[100][93]=1;ram[100][94]=1;ram[100][95]=0;ram[100][96]=1;ram[100][97]=1;ram[100][98]=1;ram[100][99]=1;ram[100][100]=0;ram[100][101]=0;ram[100][102]=1;ram[100][103]=1;ram[100][104]=1;ram[100][105]=1;ram[100][106]=0;ram[100][107]=1;ram[100][108]=1;ram[100][109]=1;ram[100][110]=1;ram[100][111]=0;ram[100][112]=1;ram[100][113]=1;ram[100][114]=1;ram[100][115]=1;ram[100][116]=1;ram[100][117]=1;ram[100][118]=1;ram[100][119]=1;ram[100][120]=1;ram[100][121]=1;ram[100][122]=1;ram[100][123]=1;ram[100][124]=0;ram[100][125]=0;ram[100][126]=1;ram[100][127]=0;ram[100][128]=0;ram[100][129]=0;ram[100][130]=0;ram[100][131]=1;ram[100][132]=1;ram[100][133]=0;ram[100][134]=1;ram[100][135]=1;ram[100][136]=1;
        ram[101][0]=1;ram[101][1]=0;ram[101][2]=1;ram[101][3]=1;ram[101][4]=1;ram[101][5]=0;ram[101][6]=1;ram[101][7]=0;ram[101][8]=1;ram[101][9]=1;ram[101][10]=1;ram[101][11]=1;ram[101][12]=0;ram[101][13]=1;ram[101][14]=1;ram[101][15]=0;ram[101][16]=1;ram[101][17]=1;ram[101][18]=1;ram[101][19]=1;ram[101][20]=1;ram[101][21]=0;ram[101][22]=1;ram[101][23]=1;ram[101][24]=1;ram[101][25]=1;ram[101][26]=1;ram[101][27]=1;ram[101][28]=1;ram[101][29]=1;ram[101][30]=1;ram[101][31]=1;ram[101][32]=1;ram[101][33]=1;ram[101][34]=1;ram[101][35]=1;ram[101][36]=1;ram[101][37]=1;ram[101][38]=0;ram[101][39]=0;ram[101][40]=1;ram[101][41]=0;ram[101][42]=1;ram[101][43]=1;ram[101][44]=1;ram[101][45]=1;ram[101][46]=0;ram[101][47]=1;ram[101][48]=1;ram[101][49]=1;ram[101][50]=1;ram[101][51]=1;ram[101][52]=0;ram[101][53]=0;ram[101][54]=1;ram[101][55]=1;ram[101][56]=1;ram[101][57]=1;ram[101][58]=1;ram[101][59]=1;ram[101][60]=1;ram[101][61]=0;ram[101][62]=1;ram[101][63]=0;ram[101][64]=1;ram[101][65]=1;ram[101][66]=1;ram[101][67]=1;ram[101][68]=0;ram[101][69]=1;ram[101][70]=0;ram[101][71]=1;ram[101][72]=0;ram[101][73]=1;ram[101][74]=1;ram[101][75]=1;ram[101][76]=1;ram[101][77]=1;ram[101][78]=0;ram[101][79]=1;ram[101][80]=1;ram[101][81]=0;ram[101][82]=1;ram[101][83]=0;ram[101][84]=1;ram[101][85]=1;ram[101][86]=1;ram[101][87]=1;ram[101][88]=1;ram[101][89]=0;ram[101][90]=0;ram[101][91]=1;ram[101][92]=1;ram[101][93]=0;ram[101][94]=1;ram[101][95]=0;ram[101][96]=1;ram[101][97]=1;ram[101][98]=1;ram[101][99]=0;ram[101][100]=0;ram[101][101]=1;ram[101][102]=1;ram[101][103]=1;ram[101][104]=1;ram[101][105]=0;ram[101][106]=1;ram[101][107]=1;ram[101][108]=1;ram[101][109]=1;ram[101][110]=0;ram[101][111]=1;ram[101][112]=0;ram[101][113]=0;ram[101][114]=1;ram[101][115]=1;ram[101][116]=0;ram[101][117]=1;ram[101][118]=1;ram[101][119]=0;ram[101][120]=1;ram[101][121]=1;ram[101][122]=1;ram[101][123]=0;ram[101][124]=1;ram[101][125]=0;ram[101][126]=1;ram[101][127]=1;ram[101][128]=0;ram[101][129]=0;ram[101][130]=1;ram[101][131]=1;ram[101][132]=1;ram[101][133]=0;ram[101][134]=0;ram[101][135]=1;ram[101][136]=1;
        ram[102][0]=0;ram[102][1]=1;ram[102][2]=1;ram[102][3]=1;ram[102][4]=1;ram[102][5]=0;ram[102][6]=1;ram[102][7]=1;ram[102][8]=0;ram[102][9]=1;ram[102][10]=1;ram[102][11]=0;ram[102][12]=1;ram[102][13]=1;ram[102][14]=1;ram[102][15]=0;ram[102][16]=1;ram[102][17]=0;ram[102][18]=1;ram[102][19]=0;ram[102][20]=1;ram[102][21]=1;ram[102][22]=1;ram[102][23]=1;ram[102][24]=1;ram[102][25]=0;ram[102][26]=1;ram[102][27]=1;ram[102][28]=1;ram[102][29]=1;ram[102][30]=0;ram[102][31]=0;ram[102][32]=1;ram[102][33]=1;ram[102][34]=1;ram[102][35]=1;ram[102][36]=1;ram[102][37]=1;ram[102][38]=0;ram[102][39]=0;ram[102][40]=1;ram[102][41]=0;ram[102][42]=1;ram[102][43]=1;ram[102][44]=1;ram[102][45]=1;ram[102][46]=0;ram[102][47]=1;ram[102][48]=1;ram[102][49]=0;ram[102][50]=1;ram[102][51]=0;ram[102][52]=1;ram[102][53]=0;ram[102][54]=1;ram[102][55]=1;ram[102][56]=0;ram[102][57]=0;ram[102][58]=1;ram[102][59]=0;ram[102][60]=0;ram[102][61]=1;ram[102][62]=1;ram[102][63]=0;ram[102][64]=0;ram[102][65]=0;ram[102][66]=0;ram[102][67]=1;ram[102][68]=1;ram[102][69]=1;ram[102][70]=1;ram[102][71]=1;ram[102][72]=0;ram[102][73]=1;ram[102][74]=0;ram[102][75]=1;ram[102][76]=0;ram[102][77]=1;ram[102][78]=1;ram[102][79]=0;ram[102][80]=0;ram[102][81]=0;ram[102][82]=1;ram[102][83]=0;ram[102][84]=1;ram[102][85]=1;ram[102][86]=1;ram[102][87]=0;ram[102][88]=0;ram[102][89]=1;ram[102][90]=1;ram[102][91]=0;ram[102][92]=1;ram[102][93]=1;ram[102][94]=1;ram[102][95]=1;ram[102][96]=1;ram[102][97]=1;ram[102][98]=1;ram[102][99]=1;ram[102][100]=0;ram[102][101]=1;ram[102][102]=0;ram[102][103]=1;ram[102][104]=1;ram[102][105]=0;ram[102][106]=0;ram[102][107]=0;ram[102][108]=1;ram[102][109]=0;ram[102][110]=1;ram[102][111]=0;ram[102][112]=0;ram[102][113]=1;ram[102][114]=1;ram[102][115]=0;ram[102][116]=1;ram[102][117]=1;ram[102][118]=1;ram[102][119]=0;ram[102][120]=1;ram[102][121]=1;ram[102][122]=1;ram[102][123]=1;ram[102][124]=1;ram[102][125]=1;ram[102][126]=1;ram[102][127]=1;ram[102][128]=1;ram[102][129]=1;ram[102][130]=1;ram[102][131]=0;ram[102][132]=1;ram[102][133]=1;ram[102][134]=0;ram[102][135]=1;ram[102][136]=1;
        ram[103][0]=1;ram[103][1]=0;ram[103][2]=1;ram[103][3]=1;ram[103][4]=0;ram[103][5]=0;ram[103][6]=0;ram[103][7]=1;ram[103][8]=1;ram[103][9]=1;ram[103][10]=0;ram[103][11]=1;ram[103][12]=1;ram[103][13]=1;ram[103][14]=0;ram[103][15]=1;ram[103][16]=1;ram[103][17]=1;ram[103][18]=1;ram[103][19]=0;ram[103][20]=1;ram[103][21]=1;ram[103][22]=1;ram[103][23]=0;ram[103][24]=0;ram[103][25]=1;ram[103][26]=1;ram[103][27]=0;ram[103][28]=1;ram[103][29]=0;ram[103][30]=1;ram[103][31]=1;ram[103][32]=1;ram[103][33]=1;ram[103][34]=1;ram[103][35]=1;ram[103][36]=1;ram[103][37]=1;ram[103][38]=1;ram[103][39]=1;ram[103][40]=0;ram[103][41]=1;ram[103][42]=1;ram[103][43]=1;ram[103][44]=1;ram[103][45]=1;ram[103][46]=0;ram[103][47]=1;ram[103][48]=1;ram[103][49]=1;ram[103][50]=1;ram[103][51]=1;ram[103][52]=1;ram[103][53]=1;ram[103][54]=0;ram[103][55]=1;ram[103][56]=0;ram[103][57]=0;ram[103][58]=0;ram[103][59]=1;ram[103][60]=1;ram[103][61]=0;ram[103][62]=1;ram[103][63]=0;ram[103][64]=1;ram[103][65]=1;ram[103][66]=1;ram[103][67]=0;ram[103][68]=1;ram[103][69]=0;ram[103][70]=1;ram[103][71]=0;ram[103][72]=1;ram[103][73]=1;ram[103][74]=1;ram[103][75]=1;ram[103][76]=0;ram[103][77]=0;ram[103][78]=1;ram[103][79]=1;ram[103][80]=0;ram[103][81]=1;ram[103][82]=1;ram[103][83]=0;ram[103][84]=1;ram[103][85]=1;ram[103][86]=0;ram[103][87]=1;ram[103][88]=1;ram[103][89]=1;ram[103][90]=1;ram[103][91]=1;ram[103][92]=0;ram[103][93]=0;ram[103][94]=1;ram[103][95]=0;ram[103][96]=1;ram[103][97]=1;ram[103][98]=1;ram[103][99]=0;ram[103][100]=0;ram[103][101]=0;ram[103][102]=0;ram[103][103]=1;ram[103][104]=1;ram[103][105]=1;ram[103][106]=1;ram[103][107]=1;ram[103][108]=1;ram[103][109]=0;ram[103][110]=0;ram[103][111]=0;ram[103][112]=0;ram[103][113]=1;ram[103][114]=1;ram[103][115]=0;ram[103][116]=0;ram[103][117]=1;ram[103][118]=0;ram[103][119]=1;ram[103][120]=1;ram[103][121]=1;ram[103][122]=1;ram[103][123]=1;ram[103][124]=1;ram[103][125]=1;ram[103][126]=1;ram[103][127]=0;ram[103][128]=0;ram[103][129]=1;ram[103][130]=1;ram[103][131]=1;ram[103][132]=1;ram[103][133]=1;ram[103][134]=1;ram[103][135]=1;ram[103][136]=1;
        ram[104][0]=0;ram[104][1]=1;ram[104][2]=0;ram[104][3]=1;ram[104][4]=1;ram[104][5]=0;ram[104][6]=1;ram[104][7]=1;ram[104][8]=0;ram[104][9]=1;ram[104][10]=0;ram[104][11]=0;ram[104][12]=1;ram[104][13]=1;ram[104][14]=1;ram[104][15]=1;ram[104][16]=1;ram[104][17]=1;ram[104][18]=1;ram[104][19]=0;ram[104][20]=1;ram[104][21]=0;ram[104][22]=1;ram[104][23]=1;ram[104][24]=1;ram[104][25]=0;ram[104][26]=0;ram[104][27]=0;ram[104][28]=1;ram[104][29]=0;ram[104][30]=1;ram[104][31]=0;ram[104][32]=1;ram[104][33]=0;ram[104][34]=1;ram[104][35]=1;ram[104][36]=1;ram[104][37]=1;ram[104][38]=1;ram[104][39]=1;ram[104][40]=1;ram[104][41]=1;ram[104][42]=0;ram[104][43]=1;ram[104][44]=1;ram[104][45]=1;ram[104][46]=0;ram[104][47]=1;ram[104][48]=1;ram[104][49]=0;ram[104][50]=1;ram[104][51]=1;ram[104][52]=1;ram[104][53]=1;ram[104][54]=1;ram[104][55]=1;ram[104][56]=1;ram[104][57]=0;ram[104][58]=1;ram[104][59]=0;ram[104][60]=1;ram[104][61]=0;ram[104][62]=1;ram[104][63]=1;ram[104][64]=1;ram[104][65]=0;ram[104][66]=1;ram[104][67]=1;ram[104][68]=1;ram[104][69]=1;ram[104][70]=1;ram[104][71]=1;ram[104][72]=1;ram[104][73]=1;ram[104][74]=0;ram[104][75]=1;ram[104][76]=0;ram[104][77]=1;ram[104][78]=1;ram[104][79]=0;ram[104][80]=0;ram[104][81]=0;ram[104][82]=1;ram[104][83]=1;ram[104][84]=0;ram[104][85]=0;ram[104][86]=1;ram[104][87]=0;ram[104][88]=0;ram[104][89]=1;ram[104][90]=1;ram[104][91]=0;ram[104][92]=1;ram[104][93]=1;ram[104][94]=1;ram[104][95]=1;ram[104][96]=0;ram[104][97]=0;ram[104][98]=1;ram[104][99]=1;ram[104][100]=0;ram[104][101]=1;ram[104][102]=1;ram[104][103]=0;ram[104][104]=1;ram[104][105]=1;ram[104][106]=1;ram[104][107]=0;ram[104][108]=0;ram[104][109]=1;ram[104][110]=0;ram[104][111]=0;ram[104][112]=1;ram[104][113]=1;ram[104][114]=0;ram[104][115]=1;ram[104][116]=1;ram[104][117]=1;ram[104][118]=0;ram[104][119]=1;ram[104][120]=1;ram[104][121]=1;ram[104][122]=1;ram[104][123]=1;ram[104][124]=1;ram[104][125]=1;ram[104][126]=1;ram[104][127]=1;ram[104][128]=1;ram[104][129]=1;ram[104][130]=0;ram[104][131]=1;ram[104][132]=0;ram[104][133]=0;ram[104][134]=1;ram[104][135]=1;ram[104][136]=1;
        ram[105][0]=1;ram[105][1]=1;ram[105][2]=1;ram[105][3]=0;ram[105][4]=0;ram[105][5]=1;ram[105][6]=1;ram[105][7]=1;ram[105][8]=1;ram[105][9]=1;ram[105][10]=1;ram[105][11]=1;ram[105][12]=1;ram[105][13]=1;ram[105][14]=1;ram[105][15]=1;ram[105][16]=1;ram[105][17]=1;ram[105][18]=0;ram[105][19]=0;ram[105][20]=1;ram[105][21]=0;ram[105][22]=1;ram[105][23]=1;ram[105][24]=1;ram[105][25]=0;ram[105][26]=0;ram[105][27]=0;ram[105][28]=1;ram[105][29]=1;ram[105][30]=0;ram[105][31]=1;ram[105][32]=1;ram[105][33]=1;ram[105][34]=1;ram[105][35]=0;ram[105][36]=0;ram[105][37]=1;ram[105][38]=1;ram[105][39]=1;ram[105][40]=1;ram[105][41]=0;ram[105][42]=1;ram[105][43]=1;ram[105][44]=0;ram[105][45]=1;ram[105][46]=1;ram[105][47]=0;ram[105][48]=1;ram[105][49]=1;ram[105][50]=1;ram[105][51]=1;ram[105][52]=1;ram[105][53]=1;ram[105][54]=0;ram[105][55]=0;ram[105][56]=0;ram[105][57]=1;ram[105][58]=0;ram[105][59]=1;ram[105][60]=0;ram[105][61]=1;ram[105][62]=1;ram[105][63]=1;ram[105][64]=1;ram[105][65]=1;ram[105][66]=0;ram[105][67]=1;ram[105][68]=0;ram[105][69]=1;ram[105][70]=1;ram[105][71]=0;ram[105][72]=1;ram[105][73]=0;ram[105][74]=1;ram[105][75]=1;ram[105][76]=1;ram[105][77]=1;ram[105][78]=1;ram[105][79]=0;ram[105][80]=1;ram[105][81]=1;ram[105][82]=1;ram[105][83]=1;ram[105][84]=0;ram[105][85]=0;ram[105][86]=0;ram[105][87]=1;ram[105][88]=0;ram[105][89]=1;ram[105][90]=1;ram[105][91]=1;ram[105][92]=0;ram[105][93]=1;ram[105][94]=0;ram[105][95]=1;ram[105][96]=1;ram[105][97]=0;ram[105][98]=1;ram[105][99]=1;ram[105][100]=1;ram[105][101]=1;ram[105][102]=1;ram[105][103]=0;ram[105][104]=1;ram[105][105]=1;ram[105][106]=1;ram[105][107]=1;ram[105][108]=0;ram[105][109]=1;ram[105][110]=0;ram[105][111]=0;ram[105][112]=1;ram[105][113]=1;ram[105][114]=1;ram[105][115]=0;ram[105][116]=0;ram[105][117]=1;ram[105][118]=0;ram[105][119]=0;ram[105][120]=1;ram[105][121]=1;ram[105][122]=1;ram[105][123]=1;ram[105][124]=0;ram[105][125]=1;ram[105][126]=1;ram[105][127]=0;ram[105][128]=1;ram[105][129]=0;ram[105][130]=0;ram[105][131]=1;ram[105][132]=0;ram[105][133]=1;ram[105][134]=1;ram[105][135]=1;ram[105][136]=0;
        ram[106][0]=1;ram[106][1]=1;ram[106][2]=1;ram[106][3]=1;ram[106][4]=0;ram[106][5]=1;ram[106][6]=1;ram[106][7]=1;ram[106][8]=0;ram[106][9]=1;ram[106][10]=0;ram[106][11]=0;ram[106][12]=0;ram[106][13]=0;ram[106][14]=1;ram[106][15]=1;ram[106][16]=1;ram[106][17]=1;ram[106][18]=1;ram[106][19]=1;ram[106][20]=1;ram[106][21]=0;ram[106][22]=1;ram[106][23]=0;ram[106][24]=0;ram[106][25]=0;ram[106][26]=0;ram[106][27]=1;ram[106][28]=1;ram[106][29]=1;ram[106][30]=0;ram[106][31]=1;ram[106][32]=0;ram[106][33]=0;ram[106][34]=0;ram[106][35]=1;ram[106][36]=1;ram[106][37]=1;ram[106][38]=1;ram[106][39]=1;ram[106][40]=0;ram[106][41]=0;ram[106][42]=0;ram[106][43]=1;ram[106][44]=1;ram[106][45]=1;ram[106][46]=1;ram[106][47]=0;ram[106][48]=1;ram[106][49]=1;ram[106][50]=0;ram[106][51]=1;ram[106][52]=1;ram[106][53]=1;ram[106][54]=1;ram[106][55]=0;ram[106][56]=0;ram[106][57]=0;ram[106][58]=0;ram[106][59]=1;ram[106][60]=0;ram[106][61]=1;ram[106][62]=1;ram[106][63]=1;ram[106][64]=1;ram[106][65]=1;ram[106][66]=0;ram[106][67]=1;ram[106][68]=1;ram[106][69]=0;ram[106][70]=1;ram[106][71]=1;ram[106][72]=1;ram[106][73]=1;ram[106][74]=1;ram[106][75]=1;ram[106][76]=1;ram[106][77]=0;ram[106][78]=0;ram[106][79]=1;ram[106][80]=1;ram[106][81]=0;ram[106][82]=1;ram[106][83]=1;ram[106][84]=0;ram[106][85]=1;ram[106][86]=0;ram[106][87]=1;ram[106][88]=1;ram[106][89]=0;ram[106][90]=1;ram[106][91]=1;ram[106][92]=1;ram[106][93]=0;ram[106][94]=1;ram[106][95]=0;ram[106][96]=1;ram[106][97]=0;ram[106][98]=1;ram[106][99]=1;ram[106][100]=0;ram[106][101]=1;ram[106][102]=0;ram[106][103]=1;ram[106][104]=1;ram[106][105]=1;ram[106][106]=1;ram[106][107]=0;ram[106][108]=1;ram[106][109]=1;ram[106][110]=0;ram[106][111]=0;ram[106][112]=1;ram[106][113]=1;ram[106][114]=1;ram[106][115]=1;ram[106][116]=0;ram[106][117]=1;ram[106][118]=1;ram[106][119]=1;ram[106][120]=1;ram[106][121]=0;ram[106][122]=1;ram[106][123]=1;ram[106][124]=1;ram[106][125]=1;ram[106][126]=1;ram[106][127]=0;ram[106][128]=0;ram[106][129]=1;ram[106][130]=0;ram[106][131]=1;ram[106][132]=0;ram[106][133]=1;ram[106][134]=0;ram[106][135]=0;ram[106][136]=1;
        ram[107][0]=1;ram[107][1]=1;ram[107][2]=0;ram[107][3]=0;ram[107][4]=1;ram[107][5]=1;ram[107][6]=1;ram[107][7]=0;ram[107][8]=0;ram[107][9]=1;ram[107][10]=1;ram[107][11]=0;ram[107][12]=1;ram[107][13]=1;ram[107][14]=1;ram[107][15]=1;ram[107][16]=0;ram[107][17]=0;ram[107][18]=0;ram[107][19]=1;ram[107][20]=0;ram[107][21]=0;ram[107][22]=1;ram[107][23]=0;ram[107][24]=0;ram[107][25]=0;ram[107][26]=0;ram[107][27]=1;ram[107][28]=0;ram[107][29]=0;ram[107][30]=0;ram[107][31]=1;ram[107][32]=0;ram[107][33]=1;ram[107][34]=0;ram[107][35]=1;ram[107][36]=1;ram[107][37]=0;ram[107][38]=1;ram[107][39]=1;ram[107][40]=1;ram[107][41]=0;ram[107][42]=1;ram[107][43]=1;ram[107][44]=1;ram[107][45]=1;ram[107][46]=1;ram[107][47]=0;ram[107][48]=0;ram[107][49]=0;ram[107][50]=0;ram[107][51]=1;ram[107][52]=1;ram[107][53]=1;ram[107][54]=1;ram[107][55]=0;ram[107][56]=1;ram[107][57]=1;ram[107][58]=0;ram[107][59]=1;ram[107][60]=0;ram[107][61]=0;ram[107][62]=1;ram[107][63]=1;ram[107][64]=1;ram[107][65]=1;ram[107][66]=0;ram[107][67]=1;ram[107][68]=1;ram[107][69]=1;ram[107][70]=1;ram[107][71]=1;ram[107][72]=0;ram[107][73]=1;ram[107][74]=1;ram[107][75]=1;ram[107][76]=0;ram[107][77]=0;ram[107][78]=1;ram[107][79]=1;ram[107][80]=1;ram[107][81]=0;ram[107][82]=1;ram[107][83]=1;ram[107][84]=0;ram[107][85]=1;ram[107][86]=0;ram[107][87]=0;ram[107][88]=1;ram[107][89]=0;ram[107][90]=0;ram[107][91]=0;ram[107][92]=1;ram[107][93]=1;ram[107][94]=1;ram[107][95]=0;ram[107][96]=1;ram[107][97]=0;ram[107][98]=0;ram[107][99]=1;ram[107][100]=1;ram[107][101]=1;ram[107][102]=0;ram[107][103]=0;ram[107][104]=1;ram[107][105]=0;ram[107][106]=1;ram[107][107]=0;ram[107][108]=1;ram[107][109]=1;ram[107][110]=0;ram[107][111]=1;ram[107][112]=0;ram[107][113]=1;ram[107][114]=0;ram[107][115]=1;ram[107][116]=0;ram[107][117]=0;ram[107][118]=0;ram[107][119]=1;ram[107][120]=1;ram[107][121]=0;ram[107][122]=1;ram[107][123]=0;ram[107][124]=1;ram[107][125]=1;ram[107][126]=1;ram[107][127]=0;ram[107][128]=1;ram[107][129]=1;ram[107][130]=0;ram[107][131]=0;ram[107][132]=1;ram[107][133]=0;ram[107][134]=1;ram[107][135]=0;ram[107][136]=0;
        ram[108][0]=0;ram[108][1]=1;ram[108][2]=0;ram[108][3]=1;ram[108][4]=0;ram[108][5]=1;ram[108][6]=0;ram[108][7]=1;ram[108][8]=1;ram[108][9]=1;ram[108][10]=1;ram[108][11]=1;ram[108][12]=0;ram[108][13]=0;ram[108][14]=1;ram[108][15]=1;ram[108][16]=1;ram[108][17]=1;ram[108][18]=1;ram[108][19]=1;ram[108][20]=0;ram[108][21]=1;ram[108][22]=1;ram[108][23]=1;ram[108][24]=1;ram[108][25]=0;ram[108][26]=1;ram[108][27]=1;ram[108][28]=1;ram[108][29]=0;ram[108][30]=0;ram[108][31]=1;ram[108][32]=1;ram[108][33]=1;ram[108][34]=1;ram[108][35]=1;ram[108][36]=1;ram[108][37]=0;ram[108][38]=1;ram[108][39]=0;ram[108][40]=0;ram[108][41]=1;ram[108][42]=0;ram[108][43]=1;ram[108][44]=1;ram[108][45]=1;ram[108][46]=1;ram[108][47]=0;ram[108][48]=0;ram[108][49]=1;ram[108][50]=1;ram[108][51]=1;ram[108][52]=1;ram[108][53]=1;ram[108][54]=0;ram[108][55]=0;ram[108][56]=1;ram[108][57]=0;ram[108][58]=1;ram[108][59]=1;ram[108][60]=1;ram[108][61]=0;ram[108][62]=0;ram[108][63]=1;ram[108][64]=1;ram[108][65]=0;ram[108][66]=1;ram[108][67]=1;ram[108][68]=0;ram[108][69]=0;ram[108][70]=0;ram[108][71]=1;ram[108][72]=1;ram[108][73]=1;ram[108][74]=1;ram[108][75]=0;ram[108][76]=1;ram[108][77]=1;ram[108][78]=1;ram[108][79]=1;ram[108][80]=0;ram[108][81]=1;ram[108][82]=1;ram[108][83]=0;ram[108][84]=1;ram[108][85]=0;ram[108][86]=1;ram[108][87]=1;ram[108][88]=0;ram[108][89]=0;ram[108][90]=1;ram[108][91]=0;ram[108][92]=0;ram[108][93]=1;ram[108][94]=1;ram[108][95]=1;ram[108][96]=0;ram[108][97]=0;ram[108][98]=1;ram[108][99]=1;ram[108][100]=1;ram[108][101]=1;ram[108][102]=0;ram[108][103]=0;ram[108][104]=1;ram[108][105]=1;ram[108][106]=1;ram[108][107]=1;ram[108][108]=1;ram[108][109]=0;ram[108][110]=0;ram[108][111]=0;ram[108][112]=1;ram[108][113]=1;ram[108][114]=0;ram[108][115]=1;ram[108][116]=1;ram[108][117]=0;ram[108][118]=0;ram[108][119]=0;ram[108][120]=1;ram[108][121]=1;ram[108][122]=0;ram[108][123]=0;ram[108][124]=1;ram[108][125]=0;ram[108][126]=1;ram[108][127]=0;ram[108][128]=0;ram[108][129]=0;ram[108][130]=0;ram[108][131]=1;ram[108][132]=1;ram[108][133]=0;ram[108][134]=1;ram[108][135]=0;ram[108][136]=1;
        ram[109][0]=1;ram[109][1]=0;ram[109][2]=0;ram[109][3]=1;ram[109][4]=1;ram[109][5]=1;ram[109][6]=0;ram[109][7]=0;ram[109][8]=0;ram[109][9]=0;ram[109][10]=0;ram[109][11]=1;ram[109][12]=0;ram[109][13]=0;ram[109][14]=1;ram[109][15]=1;ram[109][16]=1;ram[109][17]=1;ram[109][18]=0;ram[109][19]=1;ram[109][20]=0;ram[109][21]=1;ram[109][22]=1;ram[109][23]=1;ram[109][24]=1;ram[109][25]=0;ram[109][26]=1;ram[109][27]=1;ram[109][28]=1;ram[109][29]=1;ram[109][30]=0;ram[109][31]=0;ram[109][32]=1;ram[109][33]=1;ram[109][34]=1;ram[109][35]=0;ram[109][36]=1;ram[109][37]=1;ram[109][38]=1;ram[109][39]=1;ram[109][40]=0;ram[109][41]=1;ram[109][42]=0;ram[109][43]=1;ram[109][44]=1;ram[109][45]=0;ram[109][46]=0;ram[109][47]=0;ram[109][48]=1;ram[109][49]=1;ram[109][50]=1;ram[109][51]=1;ram[109][52]=0;ram[109][53]=1;ram[109][54]=1;ram[109][55]=1;ram[109][56]=1;ram[109][57]=1;ram[109][58]=1;ram[109][59]=1;ram[109][60]=1;ram[109][61]=1;ram[109][62]=0;ram[109][63]=1;ram[109][64]=0;ram[109][65]=1;ram[109][66]=1;ram[109][67]=1;ram[109][68]=0;ram[109][69]=0;ram[109][70]=0;ram[109][71]=1;ram[109][72]=1;ram[109][73]=1;ram[109][74]=0;ram[109][75]=1;ram[109][76]=0;ram[109][77]=0;ram[109][78]=1;ram[109][79]=1;ram[109][80]=0;ram[109][81]=1;ram[109][82]=0;ram[109][83]=1;ram[109][84]=0;ram[109][85]=1;ram[109][86]=1;ram[109][87]=1;ram[109][88]=1;ram[109][89]=0;ram[109][90]=0;ram[109][91]=0;ram[109][92]=1;ram[109][93]=0;ram[109][94]=1;ram[109][95]=1;ram[109][96]=1;ram[109][97]=1;ram[109][98]=0;ram[109][99]=1;ram[109][100]=1;ram[109][101]=1;ram[109][102]=1;ram[109][103]=1;ram[109][104]=0;ram[109][105]=1;ram[109][106]=1;ram[109][107]=1;ram[109][108]=1;ram[109][109]=1;ram[109][110]=1;ram[109][111]=1;ram[109][112]=1;ram[109][113]=0;ram[109][114]=1;ram[109][115]=1;ram[109][116]=0;ram[109][117]=1;ram[109][118]=1;ram[109][119]=0;ram[109][120]=1;ram[109][121]=0;ram[109][122]=1;ram[109][123]=1;ram[109][124]=1;ram[109][125]=1;ram[109][126]=1;ram[109][127]=1;ram[109][128]=1;ram[109][129]=1;ram[109][130]=1;ram[109][131]=1;ram[109][132]=0;ram[109][133]=0;ram[109][134]=0;ram[109][135]=1;ram[109][136]=1;
        ram[110][0]=1;ram[110][1]=1;ram[110][2]=1;ram[110][3]=0;ram[110][4]=1;ram[110][5]=0;ram[110][6]=1;ram[110][7]=1;ram[110][8]=1;ram[110][9]=1;ram[110][10]=1;ram[110][11]=1;ram[110][12]=1;ram[110][13]=1;ram[110][14]=1;ram[110][15]=1;ram[110][16]=1;ram[110][17]=1;ram[110][18]=1;ram[110][19]=1;ram[110][20]=0;ram[110][21]=1;ram[110][22]=1;ram[110][23]=1;ram[110][24]=0;ram[110][25]=1;ram[110][26]=1;ram[110][27]=0;ram[110][28]=0;ram[110][29]=1;ram[110][30]=1;ram[110][31]=1;ram[110][32]=1;ram[110][33]=0;ram[110][34]=1;ram[110][35]=1;ram[110][36]=1;ram[110][37]=0;ram[110][38]=1;ram[110][39]=1;ram[110][40]=0;ram[110][41]=1;ram[110][42]=0;ram[110][43]=1;ram[110][44]=1;ram[110][45]=1;ram[110][46]=1;ram[110][47]=1;ram[110][48]=1;ram[110][49]=0;ram[110][50]=0;ram[110][51]=1;ram[110][52]=1;ram[110][53]=1;ram[110][54]=1;ram[110][55]=1;ram[110][56]=1;ram[110][57]=0;ram[110][58]=1;ram[110][59]=1;ram[110][60]=0;ram[110][61]=1;ram[110][62]=1;ram[110][63]=1;ram[110][64]=1;ram[110][65]=0;ram[110][66]=1;ram[110][67]=0;ram[110][68]=0;ram[110][69]=0;ram[110][70]=1;ram[110][71]=1;ram[110][72]=0;ram[110][73]=1;ram[110][74]=1;ram[110][75]=1;ram[110][76]=1;ram[110][77]=1;ram[110][78]=0;ram[110][79]=1;ram[110][80]=1;ram[110][81]=1;ram[110][82]=1;ram[110][83]=0;ram[110][84]=0;ram[110][85]=0;ram[110][86]=1;ram[110][87]=0;ram[110][88]=0;ram[110][89]=0;ram[110][90]=1;ram[110][91]=1;ram[110][92]=0;ram[110][93]=1;ram[110][94]=1;ram[110][95]=1;ram[110][96]=1;ram[110][97]=1;ram[110][98]=0;ram[110][99]=0;ram[110][100]=1;ram[110][101]=1;ram[110][102]=1;ram[110][103]=0;ram[110][104]=1;ram[110][105]=1;ram[110][106]=0;ram[110][107]=1;ram[110][108]=1;ram[110][109]=0;ram[110][110]=0;ram[110][111]=0;ram[110][112]=1;ram[110][113]=1;ram[110][114]=1;ram[110][115]=1;ram[110][116]=1;ram[110][117]=1;ram[110][118]=1;ram[110][119]=0;ram[110][120]=0;ram[110][121]=1;ram[110][122]=1;ram[110][123]=1;ram[110][124]=1;ram[110][125]=0;ram[110][126]=0;ram[110][127]=0;ram[110][128]=1;ram[110][129]=0;ram[110][130]=0;ram[110][131]=1;ram[110][132]=1;ram[110][133]=1;ram[110][134]=0;ram[110][135]=0;ram[110][136]=1;
        ram[111][0]=1;ram[111][1]=0;ram[111][2]=1;ram[111][3]=1;ram[111][4]=1;ram[111][5]=1;ram[111][6]=0;ram[111][7]=0;ram[111][8]=1;ram[111][9]=0;ram[111][10]=0;ram[111][11]=1;ram[111][12]=1;ram[111][13]=1;ram[111][14]=1;ram[111][15]=1;ram[111][16]=1;ram[111][17]=1;ram[111][18]=1;ram[111][19]=1;ram[111][20]=0;ram[111][21]=1;ram[111][22]=1;ram[111][23]=1;ram[111][24]=1;ram[111][25]=1;ram[111][26]=0;ram[111][27]=1;ram[111][28]=1;ram[111][29]=1;ram[111][30]=1;ram[111][31]=1;ram[111][32]=0;ram[111][33]=1;ram[111][34]=1;ram[111][35]=1;ram[111][36]=1;ram[111][37]=1;ram[111][38]=0;ram[111][39]=1;ram[111][40]=1;ram[111][41]=0;ram[111][42]=1;ram[111][43]=1;ram[111][44]=0;ram[111][45]=0;ram[111][46]=1;ram[111][47]=1;ram[111][48]=0;ram[111][49]=0;ram[111][50]=0;ram[111][51]=1;ram[111][52]=1;ram[111][53]=0;ram[111][54]=1;ram[111][55]=0;ram[111][56]=0;ram[111][57]=1;ram[111][58]=1;ram[111][59]=0;ram[111][60]=1;ram[111][61]=1;ram[111][62]=1;ram[111][63]=1;ram[111][64]=1;ram[111][65]=1;ram[111][66]=1;ram[111][67]=1;ram[111][68]=0;ram[111][69]=0;ram[111][70]=0;ram[111][71]=1;ram[111][72]=1;ram[111][73]=1;ram[111][74]=0;ram[111][75]=1;ram[111][76]=1;ram[111][77]=1;ram[111][78]=1;ram[111][79]=1;ram[111][80]=1;ram[111][81]=1;ram[111][82]=1;ram[111][83]=0;ram[111][84]=0;ram[111][85]=0;ram[111][86]=1;ram[111][87]=1;ram[111][88]=1;ram[111][89]=1;ram[111][90]=1;ram[111][91]=0;ram[111][92]=0;ram[111][93]=1;ram[111][94]=1;ram[111][95]=1;ram[111][96]=0;ram[111][97]=1;ram[111][98]=0;ram[111][99]=0;ram[111][100]=1;ram[111][101]=0;ram[111][102]=1;ram[111][103]=1;ram[111][104]=1;ram[111][105]=0;ram[111][106]=1;ram[111][107]=0;ram[111][108]=0;ram[111][109]=0;ram[111][110]=1;ram[111][111]=0;ram[111][112]=1;ram[111][113]=0;ram[111][114]=1;ram[111][115]=1;ram[111][116]=1;ram[111][117]=1;ram[111][118]=1;ram[111][119]=1;ram[111][120]=1;ram[111][121]=1;ram[111][122]=1;ram[111][123]=0;ram[111][124]=1;ram[111][125]=0;ram[111][126]=0;ram[111][127]=1;ram[111][128]=1;ram[111][129]=1;ram[111][130]=1;ram[111][131]=1;ram[111][132]=1;ram[111][133]=1;ram[111][134]=1;ram[111][135]=0;ram[111][136]=1;
        ram[112][0]=1;ram[112][1]=0;ram[112][2]=1;ram[112][3]=1;ram[112][4]=1;ram[112][5]=1;ram[112][6]=1;ram[112][7]=1;ram[112][8]=1;ram[112][9]=1;ram[112][10]=0;ram[112][11]=0;ram[112][12]=1;ram[112][13]=1;ram[112][14]=1;ram[112][15]=1;ram[112][16]=0;ram[112][17]=1;ram[112][18]=1;ram[112][19]=1;ram[112][20]=1;ram[112][21]=1;ram[112][22]=1;ram[112][23]=0;ram[112][24]=0;ram[112][25]=1;ram[112][26]=1;ram[112][27]=1;ram[112][28]=0;ram[112][29]=1;ram[112][30]=1;ram[112][31]=1;ram[112][32]=0;ram[112][33]=1;ram[112][34]=1;ram[112][35]=0;ram[112][36]=0;ram[112][37]=1;ram[112][38]=1;ram[112][39]=0;ram[112][40]=1;ram[112][41]=1;ram[112][42]=1;ram[112][43]=1;ram[112][44]=1;ram[112][45]=1;ram[112][46]=1;ram[112][47]=1;ram[112][48]=1;ram[112][49]=0;ram[112][50]=1;ram[112][51]=0;ram[112][52]=1;ram[112][53]=1;ram[112][54]=0;ram[112][55]=0;ram[112][56]=0;ram[112][57]=1;ram[112][58]=1;ram[112][59]=0;ram[112][60]=0;ram[112][61]=1;ram[112][62]=1;ram[112][63]=0;ram[112][64]=1;ram[112][65]=1;ram[112][66]=1;ram[112][67]=1;ram[112][68]=0;ram[112][69]=1;ram[112][70]=1;ram[112][71]=1;ram[112][72]=1;ram[112][73]=1;ram[112][74]=1;ram[112][75]=1;ram[112][76]=1;ram[112][77]=1;ram[112][78]=1;ram[112][79]=1;ram[112][80]=1;ram[112][81]=0;ram[112][82]=1;ram[112][83]=1;ram[112][84]=1;ram[112][85]=1;ram[112][86]=1;ram[112][87]=0;ram[112][88]=1;ram[112][89]=1;ram[112][90]=0;ram[112][91]=1;ram[112][92]=0;ram[112][93]=1;ram[112][94]=1;ram[112][95]=1;ram[112][96]=0;ram[112][97]=1;ram[112][98]=0;ram[112][99]=1;ram[112][100]=1;ram[112][101]=0;ram[112][102]=0;ram[112][103]=1;ram[112][104]=1;ram[112][105]=1;ram[112][106]=1;ram[112][107]=1;ram[112][108]=1;ram[112][109]=1;ram[112][110]=1;ram[112][111]=0;ram[112][112]=1;ram[112][113]=1;ram[112][114]=0;ram[112][115]=0;ram[112][116]=1;ram[112][117]=1;ram[112][118]=1;ram[112][119]=1;ram[112][120]=1;ram[112][121]=1;ram[112][122]=1;ram[112][123]=1;ram[112][124]=0;ram[112][125]=0;ram[112][126]=1;ram[112][127]=0;ram[112][128]=0;ram[112][129]=1;ram[112][130]=1;ram[112][131]=1;ram[112][132]=1;ram[112][133]=1;ram[112][134]=1;ram[112][135]=0;ram[112][136]=0;
        ram[113][0]=1;ram[113][1]=0;ram[113][2]=1;ram[113][3]=0;ram[113][4]=1;ram[113][5]=1;ram[113][6]=0;ram[113][7]=1;ram[113][8]=1;ram[113][9]=1;ram[113][10]=1;ram[113][11]=1;ram[113][12]=0;ram[113][13]=0;ram[113][14]=0;ram[113][15]=1;ram[113][16]=1;ram[113][17]=1;ram[113][18]=0;ram[113][19]=1;ram[113][20]=0;ram[113][21]=0;ram[113][22]=1;ram[113][23]=1;ram[113][24]=1;ram[113][25]=1;ram[113][26]=0;ram[113][27]=0;ram[113][28]=1;ram[113][29]=0;ram[113][30]=0;ram[113][31]=0;ram[113][32]=1;ram[113][33]=0;ram[113][34]=0;ram[113][35]=1;ram[113][36]=1;ram[113][37]=1;ram[113][38]=1;ram[113][39]=0;ram[113][40]=0;ram[113][41]=1;ram[113][42]=0;ram[113][43]=1;ram[113][44]=0;ram[113][45]=1;ram[113][46]=1;ram[113][47]=1;ram[113][48]=0;ram[113][49]=1;ram[113][50]=1;ram[113][51]=1;ram[113][52]=1;ram[113][53]=1;ram[113][54]=1;ram[113][55]=0;ram[113][56]=1;ram[113][57]=0;ram[113][58]=0;ram[113][59]=1;ram[113][60]=1;ram[113][61]=0;ram[113][62]=1;ram[113][63]=1;ram[113][64]=1;ram[113][65]=0;ram[113][66]=1;ram[113][67]=0;ram[113][68]=1;ram[113][69]=0;ram[113][70]=0;ram[113][71]=0;ram[113][72]=1;ram[113][73]=0;ram[113][74]=1;ram[113][75]=1;ram[113][76]=1;ram[113][77]=0;ram[113][78]=1;ram[113][79]=1;ram[113][80]=1;ram[113][81]=1;ram[113][82]=0;ram[113][83]=1;ram[113][84]=1;ram[113][85]=1;ram[113][86]=0;ram[113][87]=1;ram[113][88]=1;ram[113][89]=0;ram[113][90]=1;ram[113][91]=0;ram[113][92]=1;ram[113][93]=1;ram[113][94]=1;ram[113][95]=1;ram[113][96]=1;ram[113][97]=1;ram[113][98]=1;ram[113][99]=1;ram[113][100]=1;ram[113][101]=1;ram[113][102]=0;ram[113][103]=1;ram[113][104]=1;ram[113][105]=0;ram[113][106]=1;ram[113][107]=0;ram[113][108]=1;ram[113][109]=1;ram[113][110]=1;ram[113][111]=1;ram[113][112]=1;ram[113][113]=1;ram[113][114]=1;ram[113][115]=1;ram[113][116]=1;ram[113][117]=0;ram[113][118]=0;ram[113][119]=0;ram[113][120]=1;ram[113][121]=0;ram[113][122]=1;ram[113][123]=1;ram[113][124]=0;ram[113][125]=1;ram[113][126]=1;ram[113][127]=0;ram[113][128]=1;ram[113][129]=0;ram[113][130]=0;ram[113][131]=0;ram[113][132]=1;ram[113][133]=1;ram[113][134]=1;ram[113][135]=1;ram[113][136]=1;
        ram[114][0]=0;ram[114][1]=0;ram[114][2]=1;ram[114][3]=1;ram[114][4]=1;ram[114][5]=0;ram[114][6]=0;ram[114][7]=1;ram[114][8]=1;ram[114][9]=1;ram[114][10]=0;ram[114][11]=1;ram[114][12]=0;ram[114][13]=1;ram[114][14]=1;ram[114][15]=1;ram[114][16]=1;ram[114][17]=0;ram[114][18]=1;ram[114][19]=1;ram[114][20]=1;ram[114][21]=0;ram[114][22]=1;ram[114][23]=1;ram[114][24]=0;ram[114][25]=0;ram[114][26]=1;ram[114][27]=1;ram[114][28]=0;ram[114][29]=1;ram[114][30]=0;ram[114][31]=1;ram[114][32]=0;ram[114][33]=1;ram[114][34]=0;ram[114][35]=1;ram[114][36]=1;ram[114][37]=1;ram[114][38]=0;ram[114][39]=1;ram[114][40]=0;ram[114][41]=1;ram[114][42]=1;ram[114][43]=1;ram[114][44]=1;ram[114][45]=1;ram[114][46]=1;ram[114][47]=1;ram[114][48]=1;ram[114][49]=1;ram[114][50]=0;ram[114][51]=0;ram[114][52]=1;ram[114][53]=0;ram[114][54]=1;ram[114][55]=0;ram[114][56]=0;ram[114][57]=1;ram[114][58]=0;ram[114][59]=1;ram[114][60]=1;ram[114][61]=1;ram[114][62]=0;ram[114][63]=0;ram[114][64]=1;ram[114][65]=1;ram[114][66]=0;ram[114][67]=0;ram[114][68]=0;ram[114][69]=1;ram[114][70]=1;ram[114][71]=0;ram[114][72]=0;ram[114][73]=1;ram[114][74]=0;ram[114][75]=1;ram[114][76]=0;ram[114][77]=0;ram[114][78]=1;ram[114][79]=0;ram[114][80]=0;ram[114][81]=0;ram[114][82]=1;ram[114][83]=1;ram[114][84]=1;ram[114][85]=1;ram[114][86]=0;ram[114][87]=0;ram[114][88]=1;ram[114][89]=0;ram[114][90]=1;ram[114][91]=1;ram[114][92]=0;ram[114][93]=1;ram[114][94]=1;ram[114][95]=0;ram[114][96]=1;ram[114][97]=1;ram[114][98]=1;ram[114][99]=1;ram[114][100]=1;ram[114][101]=1;ram[114][102]=0;ram[114][103]=0;ram[114][104]=1;ram[114][105]=0;ram[114][106]=0;ram[114][107]=1;ram[114][108]=1;ram[114][109]=1;ram[114][110]=0;ram[114][111]=0;ram[114][112]=0;ram[114][113]=1;ram[114][114]=1;ram[114][115]=1;ram[114][116]=0;ram[114][117]=1;ram[114][118]=0;ram[114][119]=1;ram[114][120]=1;ram[114][121]=1;ram[114][122]=0;ram[114][123]=1;ram[114][124]=0;ram[114][125]=1;ram[114][126]=1;ram[114][127]=1;ram[114][128]=0;ram[114][129]=0;ram[114][130]=0;ram[114][131]=1;ram[114][132]=1;ram[114][133]=1;ram[114][134]=1;ram[114][135]=1;ram[114][136]=0;
        ram[115][0]=0;ram[115][1]=1;ram[115][2]=0;ram[115][3]=1;ram[115][4]=1;ram[115][5]=0;ram[115][6]=1;ram[115][7]=1;ram[115][8]=1;ram[115][9]=1;ram[115][10]=0;ram[115][11]=1;ram[115][12]=1;ram[115][13]=1;ram[115][14]=1;ram[115][15]=0;ram[115][16]=0;ram[115][17]=1;ram[115][18]=1;ram[115][19]=1;ram[115][20]=0;ram[115][21]=1;ram[115][22]=0;ram[115][23]=1;ram[115][24]=1;ram[115][25]=1;ram[115][26]=1;ram[115][27]=1;ram[115][28]=1;ram[115][29]=0;ram[115][30]=1;ram[115][31]=0;ram[115][32]=0;ram[115][33]=1;ram[115][34]=1;ram[115][35]=1;ram[115][36]=0;ram[115][37]=1;ram[115][38]=1;ram[115][39]=0;ram[115][40]=1;ram[115][41]=1;ram[115][42]=1;ram[115][43]=1;ram[115][44]=1;ram[115][45]=1;ram[115][46]=1;ram[115][47]=1;ram[115][48]=0;ram[115][49]=0;ram[115][50]=1;ram[115][51]=1;ram[115][52]=1;ram[115][53]=0;ram[115][54]=0;ram[115][55]=1;ram[115][56]=0;ram[115][57]=0;ram[115][58]=1;ram[115][59]=1;ram[115][60]=1;ram[115][61]=0;ram[115][62]=0;ram[115][63]=0;ram[115][64]=1;ram[115][65]=1;ram[115][66]=1;ram[115][67]=0;ram[115][68]=1;ram[115][69]=1;ram[115][70]=0;ram[115][71]=1;ram[115][72]=1;ram[115][73]=1;ram[115][74]=0;ram[115][75]=0;ram[115][76]=0;ram[115][77]=0;ram[115][78]=1;ram[115][79]=1;ram[115][80]=1;ram[115][81]=1;ram[115][82]=1;ram[115][83]=1;ram[115][84]=1;ram[115][85]=1;ram[115][86]=1;ram[115][87]=1;ram[115][88]=1;ram[115][89]=1;ram[115][90]=1;ram[115][91]=0;ram[115][92]=0;ram[115][93]=1;ram[115][94]=1;ram[115][95]=0;ram[115][96]=1;ram[115][97]=1;ram[115][98]=1;ram[115][99]=1;ram[115][100]=0;ram[115][101]=0;ram[115][102]=1;ram[115][103]=1;ram[115][104]=1;ram[115][105]=1;ram[115][106]=0;ram[115][107]=1;ram[115][108]=0;ram[115][109]=0;ram[115][110]=1;ram[115][111]=1;ram[115][112]=1;ram[115][113]=1;ram[115][114]=0;ram[115][115]=1;ram[115][116]=0;ram[115][117]=1;ram[115][118]=0;ram[115][119]=0;ram[115][120]=1;ram[115][121]=1;ram[115][122]=1;ram[115][123]=1;ram[115][124]=1;ram[115][125]=1;ram[115][126]=1;ram[115][127]=1;ram[115][128]=0;ram[115][129]=1;ram[115][130]=0;ram[115][131]=1;ram[115][132]=0;ram[115][133]=1;ram[115][134]=0;ram[115][135]=1;ram[115][136]=1;
        ram[116][0]=1;ram[116][1]=1;ram[116][2]=1;ram[116][3]=1;ram[116][4]=0;ram[116][5]=1;ram[116][6]=1;ram[116][7]=1;ram[116][8]=1;ram[116][9]=0;ram[116][10]=1;ram[116][11]=0;ram[116][12]=0;ram[116][13]=1;ram[116][14]=1;ram[116][15]=1;ram[116][16]=0;ram[116][17]=0;ram[116][18]=1;ram[116][19]=1;ram[116][20]=1;ram[116][21]=1;ram[116][22]=0;ram[116][23]=1;ram[116][24]=1;ram[116][25]=0;ram[116][26]=1;ram[116][27]=1;ram[116][28]=0;ram[116][29]=1;ram[116][30]=0;ram[116][31]=0;ram[116][32]=1;ram[116][33]=1;ram[116][34]=1;ram[116][35]=1;ram[116][36]=1;ram[116][37]=1;ram[116][38]=0;ram[116][39]=0;ram[116][40]=0;ram[116][41]=0;ram[116][42]=1;ram[116][43]=1;ram[116][44]=1;ram[116][45]=1;ram[116][46]=1;ram[116][47]=0;ram[116][48]=0;ram[116][49]=1;ram[116][50]=1;ram[116][51]=1;ram[116][52]=1;ram[116][53]=0;ram[116][54]=0;ram[116][55]=1;ram[116][56]=1;ram[116][57]=0;ram[116][58]=1;ram[116][59]=1;ram[116][60]=1;ram[116][61]=1;ram[116][62]=1;ram[116][63]=1;ram[116][64]=0;ram[116][65]=1;ram[116][66]=0;ram[116][67]=0;ram[116][68]=0;ram[116][69]=1;ram[116][70]=0;ram[116][71]=1;ram[116][72]=1;ram[116][73]=0;ram[116][74]=0;ram[116][75]=1;ram[116][76]=1;ram[116][77]=0;ram[116][78]=1;ram[116][79]=1;ram[116][80]=1;ram[116][81]=1;ram[116][82]=1;ram[116][83]=1;ram[116][84]=1;ram[116][85]=1;ram[116][86]=0;ram[116][87]=1;ram[116][88]=0;ram[116][89]=1;ram[116][90]=1;ram[116][91]=1;ram[116][92]=1;ram[116][93]=1;ram[116][94]=0;ram[116][95]=0;ram[116][96]=0;ram[116][97]=0;ram[116][98]=0;ram[116][99]=1;ram[116][100]=0;ram[116][101]=0;ram[116][102]=1;ram[116][103]=0;ram[116][104]=1;ram[116][105]=1;ram[116][106]=1;ram[116][107]=1;ram[116][108]=0;ram[116][109]=1;ram[116][110]=1;ram[116][111]=1;ram[116][112]=0;ram[116][113]=1;ram[116][114]=1;ram[116][115]=1;ram[116][116]=0;ram[116][117]=1;ram[116][118]=1;ram[116][119]=0;ram[116][120]=0;ram[116][121]=1;ram[116][122]=1;ram[116][123]=1;ram[116][124]=1;ram[116][125]=1;ram[116][126]=1;ram[116][127]=1;ram[116][128]=1;ram[116][129]=1;ram[116][130]=0;ram[116][131]=1;ram[116][132]=0;ram[116][133]=0;ram[116][134]=1;ram[116][135]=1;ram[116][136]=0;
        ram[117][0]=0;ram[117][1]=0;ram[117][2]=1;ram[117][3]=1;ram[117][4]=1;ram[117][5]=1;ram[117][6]=1;ram[117][7]=1;ram[117][8]=1;ram[117][9]=1;ram[117][10]=0;ram[117][11]=1;ram[117][12]=1;ram[117][13]=0;ram[117][14]=0;ram[117][15]=1;ram[117][16]=1;ram[117][17]=1;ram[117][18]=0;ram[117][19]=1;ram[117][20]=1;ram[117][21]=0;ram[117][22]=1;ram[117][23]=0;ram[117][24]=0;ram[117][25]=0;ram[117][26]=1;ram[117][27]=1;ram[117][28]=1;ram[117][29]=0;ram[117][30]=0;ram[117][31]=1;ram[117][32]=0;ram[117][33]=0;ram[117][34]=1;ram[117][35]=0;ram[117][36]=0;ram[117][37]=1;ram[117][38]=1;ram[117][39]=1;ram[117][40]=0;ram[117][41]=0;ram[117][42]=1;ram[117][43]=1;ram[117][44]=1;ram[117][45]=1;ram[117][46]=1;ram[117][47]=0;ram[117][48]=1;ram[117][49]=1;ram[117][50]=1;ram[117][51]=0;ram[117][52]=0;ram[117][53]=1;ram[117][54]=1;ram[117][55]=1;ram[117][56]=1;ram[117][57]=0;ram[117][58]=1;ram[117][59]=0;ram[117][60]=1;ram[117][61]=0;ram[117][62]=1;ram[117][63]=0;ram[117][64]=1;ram[117][65]=0;ram[117][66]=1;ram[117][67]=1;ram[117][68]=0;ram[117][69]=1;ram[117][70]=1;ram[117][71]=1;ram[117][72]=1;ram[117][73]=1;ram[117][74]=1;ram[117][75]=0;ram[117][76]=1;ram[117][77]=1;ram[117][78]=0;ram[117][79]=1;ram[117][80]=1;ram[117][81]=0;ram[117][82]=1;ram[117][83]=1;ram[117][84]=1;ram[117][85]=1;ram[117][86]=0;ram[117][87]=1;ram[117][88]=1;ram[117][89]=0;ram[117][90]=0;ram[117][91]=0;ram[117][92]=1;ram[117][93]=0;ram[117][94]=1;ram[117][95]=1;ram[117][96]=1;ram[117][97]=1;ram[117][98]=1;ram[117][99]=1;ram[117][100]=0;ram[117][101]=1;ram[117][102]=0;ram[117][103]=1;ram[117][104]=0;ram[117][105]=1;ram[117][106]=1;ram[117][107]=1;ram[117][108]=0;ram[117][109]=0;ram[117][110]=0;ram[117][111]=1;ram[117][112]=1;ram[117][113]=1;ram[117][114]=1;ram[117][115]=0;ram[117][116]=1;ram[117][117]=1;ram[117][118]=1;ram[117][119]=0;ram[117][120]=1;ram[117][121]=1;ram[117][122]=1;ram[117][123]=0;ram[117][124]=1;ram[117][125]=0;ram[117][126]=1;ram[117][127]=1;ram[117][128]=0;ram[117][129]=0;ram[117][130]=1;ram[117][131]=1;ram[117][132]=1;ram[117][133]=1;ram[117][134]=0;ram[117][135]=0;ram[117][136]=1;
        ram[118][0]=0;ram[118][1]=0;ram[118][2]=1;ram[118][3]=1;ram[118][4]=0;ram[118][5]=1;ram[118][6]=0;ram[118][7]=0;ram[118][8]=1;ram[118][9]=1;ram[118][10]=1;ram[118][11]=1;ram[118][12]=1;ram[118][13]=1;ram[118][14]=1;ram[118][15]=1;ram[118][16]=1;ram[118][17]=1;ram[118][18]=1;ram[118][19]=1;ram[118][20]=1;ram[118][21]=1;ram[118][22]=0;ram[118][23]=1;ram[118][24]=1;ram[118][25]=1;ram[118][26]=1;ram[118][27]=0;ram[118][28]=1;ram[118][29]=1;ram[118][30]=1;ram[118][31]=0;ram[118][32]=1;ram[118][33]=1;ram[118][34]=1;ram[118][35]=1;ram[118][36]=1;ram[118][37]=1;ram[118][38]=0;ram[118][39]=1;ram[118][40]=1;ram[118][41]=1;ram[118][42]=1;ram[118][43]=1;ram[118][44]=0;ram[118][45]=0;ram[118][46]=1;ram[118][47]=1;ram[118][48]=0;ram[118][49]=0;ram[118][50]=0;ram[118][51]=1;ram[118][52]=1;ram[118][53]=0;ram[118][54]=0;ram[118][55]=0;ram[118][56]=1;ram[118][57]=1;ram[118][58]=1;ram[118][59]=0;ram[118][60]=1;ram[118][61]=0;ram[118][62]=0;ram[118][63]=1;ram[118][64]=1;ram[118][65]=0;ram[118][66]=1;ram[118][67]=0;ram[118][68]=1;ram[118][69]=1;ram[118][70]=0;ram[118][71]=1;ram[118][72]=0;ram[118][73]=0;ram[118][74]=0;ram[118][75]=1;ram[118][76]=0;ram[118][77]=1;ram[118][78]=1;ram[118][79]=0;ram[118][80]=1;ram[118][81]=1;ram[118][82]=0;ram[118][83]=0;ram[118][84]=1;ram[118][85]=1;ram[118][86]=1;ram[118][87]=1;ram[118][88]=0;ram[118][89]=1;ram[118][90]=0;ram[118][91]=0;ram[118][92]=1;ram[118][93]=1;ram[118][94]=1;ram[118][95]=0;ram[118][96]=0;ram[118][97]=0;ram[118][98]=0;ram[118][99]=1;ram[118][100]=0;ram[118][101]=1;ram[118][102]=1;ram[118][103]=1;ram[118][104]=1;ram[118][105]=0;ram[118][106]=1;ram[118][107]=0;ram[118][108]=0;ram[118][109]=0;ram[118][110]=1;ram[118][111]=1;ram[118][112]=1;ram[118][113]=1;ram[118][114]=0;ram[118][115]=1;ram[118][116]=1;ram[118][117]=1;ram[118][118]=0;ram[118][119]=0;ram[118][120]=1;ram[118][121]=1;ram[118][122]=0;ram[118][123]=0;ram[118][124]=1;ram[118][125]=1;ram[118][126]=1;ram[118][127]=1;ram[118][128]=1;ram[118][129]=0;ram[118][130]=1;ram[118][131]=1;ram[118][132]=1;ram[118][133]=1;ram[118][134]=1;ram[118][135]=1;ram[118][136]=1;
        ram[119][0]=1;ram[119][1]=1;ram[119][2]=1;ram[119][3]=1;ram[119][4]=1;ram[119][5]=0;ram[119][6]=1;ram[119][7]=1;ram[119][8]=1;ram[119][9]=0;ram[119][10]=0;ram[119][11]=1;ram[119][12]=1;ram[119][13]=0;ram[119][14]=0;ram[119][15]=1;ram[119][16]=0;ram[119][17]=1;ram[119][18]=0;ram[119][19]=0;ram[119][20]=0;ram[119][21]=1;ram[119][22]=0;ram[119][23]=0;ram[119][24]=1;ram[119][25]=1;ram[119][26]=0;ram[119][27]=0;ram[119][28]=0;ram[119][29]=0;ram[119][30]=0;ram[119][31]=1;ram[119][32]=0;ram[119][33]=1;ram[119][34]=0;ram[119][35]=1;ram[119][36]=1;ram[119][37]=0;ram[119][38]=0;ram[119][39]=0;ram[119][40]=1;ram[119][41]=0;ram[119][42]=1;ram[119][43]=0;ram[119][44]=1;ram[119][45]=0;ram[119][46]=1;ram[119][47]=1;ram[119][48]=0;ram[119][49]=1;ram[119][50]=0;ram[119][51]=1;ram[119][52]=1;ram[119][53]=0;ram[119][54]=0;ram[119][55]=1;ram[119][56]=1;ram[119][57]=1;ram[119][58]=1;ram[119][59]=0;ram[119][60]=0;ram[119][61]=1;ram[119][62]=1;ram[119][63]=1;ram[119][64]=1;ram[119][65]=1;ram[119][66]=1;ram[119][67]=1;ram[119][68]=1;ram[119][69]=0;ram[119][70]=1;ram[119][71]=0;ram[119][72]=1;ram[119][73]=1;ram[119][74]=1;ram[119][75]=1;ram[119][76]=1;ram[119][77]=1;ram[119][78]=0;ram[119][79]=1;ram[119][80]=1;ram[119][81]=1;ram[119][82]=0;ram[119][83]=1;ram[119][84]=1;ram[119][85]=1;ram[119][86]=1;ram[119][87]=1;ram[119][88]=0;ram[119][89]=0;ram[119][90]=0;ram[119][91]=1;ram[119][92]=1;ram[119][93]=0;ram[119][94]=1;ram[119][95]=0;ram[119][96]=1;ram[119][97]=1;ram[119][98]=1;ram[119][99]=0;ram[119][100]=0;ram[119][101]=1;ram[119][102]=1;ram[119][103]=1;ram[119][104]=1;ram[119][105]=0;ram[119][106]=1;ram[119][107]=1;ram[119][108]=1;ram[119][109]=0;ram[119][110]=1;ram[119][111]=1;ram[119][112]=0;ram[119][113]=1;ram[119][114]=1;ram[119][115]=0;ram[119][116]=1;ram[119][117]=1;ram[119][118]=0;ram[119][119]=1;ram[119][120]=1;ram[119][121]=0;ram[119][122]=1;ram[119][123]=1;ram[119][124]=1;ram[119][125]=1;ram[119][126]=1;ram[119][127]=1;ram[119][128]=0;ram[119][129]=0;ram[119][130]=1;ram[119][131]=1;ram[119][132]=0;ram[119][133]=1;ram[119][134]=0;ram[119][135]=1;ram[119][136]=1;
        ram[120][0]=1;ram[120][1]=1;ram[120][2]=1;ram[120][3]=1;ram[120][4]=1;ram[120][5]=1;ram[120][6]=1;ram[120][7]=1;ram[120][8]=0;ram[120][9]=0;ram[120][10]=1;ram[120][11]=1;ram[120][12]=1;ram[120][13]=1;ram[120][14]=1;ram[120][15]=1;ram[120][16]=0;ram[120][17]=1;ram[120][18]=0;ram[120][19]=0;ram[120][20]=1;ram[120][21]=0;ram[120][22]=1;ram[120][23]=0;ram[120][24]=1;ram[120][25]=0;ram[120][26]=1;ram[120][27]=1;ram[120][28]=1;ram[120][29]=1;ram[120][30]=1;ram[120][31]=1;ram[120][32]=1;ram[120][33]=0;ram[120][34]=0;ram[120][35]=1;ram[120][36]=0;ram[120][37]=1;ram[120][38]=1;ram[120][39]=1;ram[120][40]=1;ram[120][41]=1;ram[120][42]=0;ram[120][43]=1;ram[120][44]=0;ram[120][45]=0;ram[120][46]=1;ram[120][47]=1;ram[120][48]=1;ram[120][49]=0;ram[120][50]=1;ram[120][51]=1;ram[120][52]=1;ram[120][53]=1;ram[120][54]=1;ram[120][55]=1;ram[120][56]=1;ram[120][57]=1;ram[120][58]=1;ram[120][59]=1;ram[120][60]=1;ram[120][61]=1;ram[120][62]=1;ram[120][63]=0;ram[120][64]=1;ram[120][65]=1;ram[120][66]=0;ram[120][67]=0;ram[120][68]=1;ram[120][69]=0;ram[120][70]=0;ram[120][71]=1;ram[120][72]=0;ram[120][73]=1;ram[120][74]=1;ram[120][75]=1;ram[120][76]=1;ram[120][77]=1;ram[120][78]=1;ram[120][79]=1;ram[120][80]=0;ram[120][81]=1;ram[120][82]=0;ram[120][83]=1;ram[120][84]=0;ram[120][85]=1;ram[120][86]=0;ram[120][87]=1;ram[120][88]=1;ram[120][89]=1;ram[120][90]=0;ram[120][91]=1;ram[120][92]=0;ram[120][93]=0;ram[120][94]=1;ram[120][95]=1;ram[120][96]=1;ram[120][97]=1;ram[120][98]=1;ram[120][99]=1;ram[120][100]=1;ram[120][101]=0;ram[120][102]=0;ram[120][103]=1;ram[120][104]=1;ram[120][105]=1;ram[120][106]=1;ram[120][107]=0;ram[120][108]=0;ram[120][109]=1;ram[120][110]=1;ram[120][111]=1;ram[120][112]=1;ram[120][113]=1;ram[120][114]=0;ram[120][115]=1;ram[120][116]=1;ram[120][117]=1;ram[120][118]=0;ram[120][119]=1;ram[120][120]=1;ram[120][121]=1;ram[120][122]=0;ram[120][123]=1;ram[120][124]=1;ram[120][125]=1;ram[120][126]=1;ram[120][127]=1;ram[120][128]=1;ram[120][129]=1;ram[120][130]=1;ram[120][131]=1;ram[120][132]=0;ram[120][133]=0;ram[120][134]=0;ram[120][135]=1;ram[120][136]=1;
        ram[121][0]=0;ram[121][1]=0;ram[121][2]=1;ram[121][3]=1;ram[121][4]=0;ram[121][5]=1;ram[121][6]=1;ram[121][7]=0;ram[121][8]=0;ram[121][9]=1;ram[121][10]=1;ram[121][11]=1;ram[121][12]=0;ram[121][13]=1;ram[121][14]=1;ram[121][15]=1;ram[121][16]=1;ram[121][17]=1;ram[121][18]=1;ram[121][19]=1;ram[121][20]=0;ram[121][21]=1;ram[121][22]=1;ram[121][23]=0;ram[121][24]=1;ram[121][25]=1;ram[121][26]=1;ram[121][27]=1;ram[121][28]=1;ram[121][29]=0;ram[121][30]=1;ram[121][31]=0;ram[121][32]=1;ram[121][33]=1;ram[121][34]=0;ram[121][35]=0;ram[121][36]=1;ram[121][37]=0;ram[121][38]=1;ram[121][39]=1;ram[121][40]=1;ram[121][41]=1;ram[121][42]=1;ram[121][43]=1;ram[121][44]=1;ram[121][45]=0;ram[121][46]=1;ram[121][47]=0;ram[121][48]=0;ram[121][49]=1;ram[121][50]=1;ram[121][51]=1;ram[121][52]=1;ram[121][53]=1;ram[121][54]=0;ram[121][55]=0;ram[121][56]=0;ram[121][57]=1;ram[121][58]=1;ram[121][59]=1;ram[121][60]=1;ram[121][61]=1;ram[121][62]=0;ram[121][63]=0;ram[121][64]=0;ram[121][65]=1;ram[121][66]=1;ram[121][67]=1;ram[121][68]=1;ram[121][69]=1;ram[121][70]=1;ram[121][71]=1;ram[121][72]=0;ram[121][73]=0;ram[121][74]=1;ram[121][75]=1;ram[121][76]=1;ram[121][77]=1;ram[121][78]=1;ram[121][79]=1;ram[121][80]=1;ram[121][81]=1;ram[121][82]=1;ram[121][83]=0;ram[121][84]=1;ram[121][85]=1;ram[121][86]=1;ram[121][87]=1;ram[121][88]=0;ram[121][89]=1;ram[121][90]=1;ram[121][91]=1;ram[121][92]=1;ram[121][93]=1;ram[121][94]=1;ram[121][95]=0;ram[121][96]=1;ram[121][97]=1;ram[121][98]=0;ram[121][99]=0;ram[121][100]=1;ram[121][101]=0;ram[121][102]=1;ram[121][103]=1;ram[121][104]=1;ram[121][105]=1;ram[121][106]=1;ram[121][107]=1;ram[121][108]=1;ram[121][109]=1;ram[121][110]=1;ram[121][111]=1;ram[121][112]=1;ram[121][113]=1;ram[121][114]=1;ram[121][115]=1;ram[121][116]=1;ram[121][117]=0;ram[121][118]=1;ram[121][119]=1;ram[121][120]=1;ram[121][121]=0;ram[121][122]=1;ram[121][123]=1;ram[121][124]=0;ram[121][125]=1;ram[121][126]=0;ram[121][127]=0;ram[121][128]=1;ram[121][129]=1;ram[121][130]=1;ram[121][131]=1;ram[121][132]=1;ram[121][133]=1;ram[121][134]=1;ram[121][135]=1;ram[121][136]=1;
        ram[122][0]=0;ram[122][1]=0;ram[122][2]=1;ram[122][3]=1;ram[122][4]=1;ram[122][5]=1;ram[122][6]=0;ram[122][7]=1;ram[122][8]=1;ram[122][9]=1;ram[122][10]=1;ram[122][11]=0;ram[122][12]=1;ram[122][13]=1;ram[122][14]=1;ram[122][15]=0;ram[122][16]=0;ram[122][17]=1;ram[122][18]=1;ram[122][19]=1;ram[122][20]=0;ram[122][21]=1;ram[122][22]=1;ram[122][23]=0;ram[122][24]=0;ram[122][25]=1;ram[122][26]=1;ram[122][27]=1;ram[122][28]=1;ram[122][29]=1;ram[122][30]=1;ram[122][31]=0;ram[122][32]=1;ram[122][33]=1;ram[122][34]=0;ram[122][35]=1;ram[122][36]=0;ram[122][37]=0;ram[122][38]=0;ram[122][39]=1;ram[122][40]=0;ram[122][41]=0;ram[122][42]=1;ram[122][43]=1;ram[122][44]=1;ram[122][45]=1;ram[122][46]=0;ram[122][47]=1;ram[122][48]=0;ram[122][49]=1;ram[122][50]=1;ram[122][51]=1;ram[122][52]=0;ram[122][53]=1;ram[122][54]=1;ram[122][55]=1;ram[122][56]=1;ram[122][57]=1;ram[122][58]=0;ram[122][59]=1;ram[122][60]=1;ram[122][61]=0;ram[122][62]=0;ram[122][63]=1;ram[122][64]=1;ram[122][65]=1;ram[122][66]=0;ram[122][67]=1;ram[122][68]=1;ram[122][69]=0;ram[122][70]=0;ram[122][71]=1;ram[122][72]=1;ram[122][73]=1;ram[122][74]=1;ram[122][75]=0;ram[122][76]=1;ram[122][77]=0;ram[122][78]=0;ram[122][79]=0;ram[122][80]=1;ram[122][81]=1;ram[122][82]=1;ram[122][83]=0;ram[122][84]=1;ram[122][85]=1;ram[122][86]=1;ram[122][87]=0;ram[122][88]=1;ram[122][89]=1;ram[122][90]=1;ram[122][91]=1;ram[122][92]=1;ram[122][93]=1;ram[122][94]=1;ram[122][95]=1;ram[122][96]=1;ram[122][97]=1;ram[122][98]=1;ram[122][99]=0;ram[122][100]=1;ram[122][101]=1;ram[122][102]=1;ram[122][103]=0;ram[122][104]=0;ram[122][105]=1;ram[122][106]=0;ram[122][107]=0;ram[122][108]=1;ram[122][109]=1;ram[122][110]=1;ram[122][111]=1;ram[122][112]=0;ram[122][113]=1;ram[122][114]=1;ram[122][115]=1;ram[122][116]=1;ram[122][117]=0;ram[122][118]=1;ram[122][119]=1;ram[122][120]=1;ram[122][121]=0;ram[122][122]=0;ram[122][123]=1;ram[122][124]=1;ram[122][125]=1;ram[122][126]=0;ram[122][127]=0;ram[122][128]=0;ram[122][129]=1;ram[122][130]=0;ram[122][131]=1;ram[122][132]=1;ram[122][133]=0;ram[122][134]=1;ram[122][135]=1;ram[122][136]=1;
        ram[123][0]=1;ram[123][1]=1;ram[123][2]=1;ram[123][3]=1;ram[123][4]=0;ram[123][5]=1;ram[123][6]=0;ram[123][7]=0;ram[123][8]=0;ram[123][9]=1;ram[123][10]=0;ram[123][11]=1;ram[123][12]=1;ram[123][13]=1;ram[123][14]=0;ram[123][15]=0;ram[123][16]=1;ram[123][17]=1;ram[123][18]=1;ram[123][19]=1;ram[123][20]=1;ram[123][21]=0;ram[123][22]=1;ram[123][23]=1;ram[123][24]=1;ram[123][25]=0;ram[123][26]=1;ram[123][27]=0;ram[123][28]=1;ram[123][29]=1;ram[123][30]=1;ram[123][31]=0;ram[123][32]=1;ram[123][33]=0;ram[123][34]=1;ram[123][35]=0;ram[123][36]=1;ram[123][37]=1;ram[123][38]=0;ram[123][39]=1;ram[123][40]=1;ram[123][41]=0;ram[123][42]=1;ram[123][43]=1;ram[123][44]=1;ram[123][45]=0;ram[123][46]=1;ram[123][47]=1;ram[123][48]=1;ram[123][49]=0;ram[123][50]=0;ram[123][51]=1;ram[123][52]=1;ram[123][53]=1;ram[123][54]=1;ram[123][55]=0;ram[123][56]=0;ram[123][57]=1;ram[123][58]=1;ram[123][59]=0;ram[123][60]=1;ram[123][61]=1;ram[123][62]=1;ram[123][63]=1;ram[123][64]=1;ram[123][65]=1;ram[123][66]=1;ram[123][67]=0;ram[123][68]=1;ram[123][69]=0;ram[123][70]=1;ram[123][71]=1;ram[123][72]=0;ram[123][73]=0;ram[123][74]=0;ram[123][75]=0;ram[123][76]=0;ram[123][77]=0;ram[123][78]=1;ram[123][79]=0;ram[123][80]=1;ram[123][81]=1;ram[123][82]=0;ram[123][83]=1;ram[123][84]=1;ram[123][85]=1;ram[123][86]=0;ram[123][87]=1;ram[123][88]=0;ram[123][89]=1;ram[123][90]=1;ram[123][91]=0;ram[123][92]=0;ram[123][93]=1;ram[123][94]=1;ram[123][95]=1;ram[123][96]=1;ram[123][97]=1;ram[123][98]=1;ram[123][99]=1;ram[123][100]=1;ram[123][101]=1;ram[123][102]=0;ram[123][103]=0;ram[123][104]=0;ram[123][105]=1;ram[123][106]=1;ram[123][107]=1;ram[123][108]=0;ram[123][109]=1;ram[123][110]=1;ram[123][111]=0;ram[123][112]=0;ram[123][113]=1;ram[123][114]=1;ram[123][115]=0;ram[123][116]=0;ram[123][117]=1;ram[123][118]=1;ram[123][119]=1;ram[123][120]=1;ram[123][121]=0;ram[123][122]=1;ram[123][123]=1;ram[123][124]=1;ram[123][125]=1;ram[123][126]=0;ram[123][127]=1;ram[123][128]=1;ram[123][129]=1;ram[123][130]=1;ram[123][131]=0;ram[123][132]=0;ram[123][133]=1;ram[123][134]=1;ram[123][135]=1;ram[123][136]=1;
        ram[124][0]=1;ram[124][1]=0;ram[124][2]=0;ram[124][3]=1;ram[124][4]=1;ram[124][5]=1;ram[124][6]=1;ram[124][7]=1;ram[124][8]=1;ram[124][9]=1;ram[124][10]=1;ram[124][11]=1;ram[124][12]=0;ram[124][13]=0;ram[124][14]=1;ram[124][15]=0;ram[124][16]=0;ram[124][17]=0;ram[124][18]=1;ram[124][19]=1;ram[124][20]=1;ram[124][21]=1;ram[124][22]=0;ram[124][23]=1;ram[124][24]=1;ram[124][25]=0;ram[124][26]=0;ram[124][27]=0;ram[124][28]=0;ram[124][29]=1;ram[124][30]=1;ram[124][31]=1;ram[124][32]=1;ram[124][33]=1;ram[124][34]=1;ram[124][35]=0;ram[124][36]=0;ram[124][37]=1;ram[124][38]=1;ram[124][39]=1;ram[124][40]=1;ram[124][41]=1;ram[124][42]=1;ram[124][43]=1;ram[124][44]=0;ram[124][45]=1;ram[124][46]=1;ram[124][47]=0;ram[124][48]=1;ram[124][49]=1;ram[124][50]=1;ram[124][51]=0;ram[124][52]=0;ram[124][53]=1;ram[124][54]=0;ram[124][55]=0;ram[124][56]=1;ram[124][57]=0;ram[124][58]=0;ram[124][59]=0;ram[124][60]=1;ram[124][61]=1;ram[124][62]=1;ram[124][63]=1;ram[124][64]=0;ram[124][65]=1;ram[124][66]=0;ram[124][67]=1;ram[124][68]=1;ram[124][69]=1;ram[124][70]=1;ram[124][71]=0;ram[124][72]=1;ram[124][73]=0;ram[124][74]=0;ram[124][75]=1;ram[124][76]=0;ram[124][77]=1;ram[124][78]=1;ram[124][79]=0;ram[124][80]=1;ram[124][81]=1;ram[124][82]=0;ram[124][83]=1;ram[124][84]=1;ram[124][85]=1;ram[124][86]=1;ram[124][87]=1;ram[124][88]=1;ram[124][89]=1;ram[124][90]=1;ram[124][91]=1;ram[124][92]=1;ram[124][93]=1;ram[124][94]=0;ram[124][95]=1;ram[124][96]=0;ram[124][97]=0;ram[124][98]=1;ram[124][99]=0;ram[124][100]=0;ram[124][101]=1;ram[124][102]=1;ram[124][103]=0;ram[124][104]=0;ram[124][105]=0;ram[124][106]=1;ram[124][107]=0;ram[124][108]=1;ram[124][109]=0;ram[124][110]=1;ram[124][111]=0;ram[124][112]=1;ram[124][113]=1;ram[124][114]=0;ram[124][115]=0;ram[124][116]=1;ram[124][117]=1;ram[124][118]=1;ram[124][119]=1;ram[124][120]=1;ram[124][121]=1;ram[124][122]=0;ram[124][123]=1;ram[124][124]=0;ram[124][125]=1;ram[124][126]=0;ram[124][127]=1;ram[124][128]=1;ram[124][129]=0;ram[124][130]=0;ram[124][131]=0;ram[124][132]=1;ram[124][133]=1;ram[124][134]=1;ram[124][135]=1;ram[124][136]=1;
        ram[125][0]=0;ram[125][1]=1;ram[125][2]=1;ram[125][3]=1;ram[125][4]=1;ram[125][5]=0;ram[125][6]=0;ram[125][7]=1;ram[125][8]=1;ram[125][9]=1;ram[125][10]=1;ram[125][11]=1;ram[125][12]=1;ram[125][13]=1;ram[125][14]=1;ram[125][15]=0;ram[125][16]=1;ram[125][17]=0;ram[125][18]=0;ram[125][19]=1;ram[125][20]=1;ram[125][21]=0;ram[125][22]=1;ram[125][23]=1;ram[125][24]=1;ram[125][25]=1;ram[125][26]=0;ram[125][27]=1;ram[125][28]=1;ram[125][29]=1;ram[125][30]=1;ram[125][31]=1;ram[125][32]=0;ram[125][33]=0;ram[125][34]=0;ram[125][35]=0;ram[125][36]=1;ram[125][37]=0;ram[125][38]=1;ram[125][39]=0;ram[125][40]=1;ram[125][41]=0;ram[125][42]=1;ram[125][43]=0;ram[125][44]=1;ram[125][45]=1;ram[125][46]=0;ram[125][47]=1;ram[125][48]=0;ram[125][49]=1;ram[125][50]=0;ram[125][51]=0;ram[125][52]=0;ram[125][53]=1;ram[125][54]=1;ram[125][55]=0;ram[125][56]=0;ram[125][57]=1;ram[125][58]=1;ram[125][59]=0;ram[125][60]=1;ram[125][61]=1;ram[125][62]=1;ram[125][63]=0;ram[125][64]=1;ram[125][65]=1;ram[125][66]=0;ram[125][67]=1;ram[125][68]=1;ram[125][69]=0;ram[125][70]=0;ram[125][71]=1;ram[125][72]=0;ram[125][73]=1;ram[125][74]=1;ram[125][75]=1;ram[125][76]=1;ram[125][77]=1;ram[125][78]=0;ram[125][79]=0;ram[125][80]=1;ram[125][81]=0;ram[125][82]=0;ram[125][83]=1;ram[125][84]=1;ram[125][85]=1;ram[125][86]=0;ram[125][87]=0;ram[125][88]=1;ram[125][89]=1;ram[125][90]=1;ram[125][91]=0;ram[125][92]=1;ram[125][93]=0;ram[125][94]=1;ram[125][95]=0;ram[125][96]=1;ram[125][97]=0;ram[125][98]=1;ram[125][99]=1;ram[125][100]=1;ram[125][101]=1;ram[125][102]=1;ram[125][103]=0;ram[125][104]=0;ram[125][105]=1;ram[125][106]=0;ram[125][107]=1;ram[125][108]=0;ram[125][109]=0;ram[125][110]=1;ram[125][111]=1;ram[125][112]=0;ram[125][113]=0;ram[125][114]=1;ram[125][115]=1;ram[125][116]=1;ram[125][117]=1;ram[125][118]=0;ram[125][119]=1;ram[125][120]=0;ram[125][121]=1;ram[125][122]=1;ram[125][123]=1;ram[125][124]=0;ram[125][125]=1;ram[125][126]=1;ram[125][127]=0;ram[125][128]=1;ram[125][129]=1;ram[125][130]=0;ram[125][131]=0;ram[125][132]=0;ram[125][133]=0;ram[125][134]=1;ram[125][135]=1;ram[125][136]=0;
        ram[126][0]=1;ram[126][1]=1;ram[126][2]=0;ram[126][3]=1;ram[126][4]=1;ram[126][5]=1;ram[126][6]=1;ram[126][7]=1;ram[126][8]=1;ram[126][9]=0;ram[126][10]=0;ram[126][11]=1;ram[126][12]=0;ram[126][13]=0;ram[126][14]=0;ram[126][15]=1;ram[126][16]=1;ram[126][17]=1;ram[126][18]=1;ram[126][19]=0;ram[126][20]=1;ram[126][21]=1;ram[126][22]=1;ram[126][23]=0;ram[126][24]=0;ram[126][25]=1;ram[126][26]=0;ram[126][27]=1;ram[126][28]=1;ram[126][29]=0;ram[126][30]=0;ram[126][31]=0;ram[126][32]=0;ram[126][33]=1;ram[126][34]=1;ram[126][35]=0;ram[126][36]=0;ram[126][37]=1;ram[126][38]=1;ram[126][39]=1;ram[126][40]=1;ram[126][41]=1;ram[126][42]=1;ram[126][43]=0;ram[126][44]=0;ram[126][45]=0;ram[126][46]=0;ram[126][47]=0;ram[126][48]=1;ram[126][49]=1;ram[126][50]=0;ram[126][51]=1;ram[126][52]=1;ram[126][53]=1;ram[126][54]=1;ram[126][55]=1;ram[126][56]=1;ram[126][57]=1;ram[126][58]=0;ram[126][59]=0;ram[126][60]=1;ram[126][61]=1;ram[126][62]=1;ram[126][63]=0;ram[126][64]=0;ram[126][65]=1;ram[126][66]=1;ram[126][67]=0;ram[126][68]=1;ram[126][69]=1;ram[126][70]=1;ram[126][71]=1;ram[126][72]=1;ram[126][73]=1;ram[126][74]=1;ram[126][75]=1;ram[126][76]=0;ram[126][77]=0;ram[126][78]=1;ram[126][79]=1;ram[126][80]=1;ram[126][81]=1;ram[126][82]=0;ram[126][83]=1;ram[126][84]=0;ram[126][85]=0;ram[126][86]=0;ram[126][87]=1;ram[126][88]=0;ram[126][89]=1;ram[126][90]=1;ram[126][91]=1;ram[126][92]=1;ram[126][93]=1;ram[126][94]=0;ram[126][95]=1;ram[126][96]=0;ram[126][97]=1;ram[126][98]=1;ram[126][99]=1;ram[126][100]=1;ram[126][101]=0;ram[126][102]=1;ram[126][103]=0;ram[126][104]=1;ram[126][105]=1;ram[126][106]=1;ram[126][107]=1;ram[126][108]=0;ram[126][109]=1;ram[126][110]=0;ram[126][111]=0;ram[126][112]=1;ram[126][113]=0;ram[126][114]=0;ram[126][115]=1;ram[126][116]=1;ram[126][117]=1;ram[126][118]=1;ram[126][119]=1;ram[126][120]=0;ram[126][121]=1;ram[126][122]=1;ram[126][123]=1;ram[126][124]=0;ram[126][125]=0;ram[126][126]=0;ram[126][127]=0;ram[126][128]=1;ram[126][129]=0;ram[126][130]=1;ram[126][131]=1;ram[126][132]=1;ram[126][133]=0;ram[126][134]=1;ram[126][135]=1;ram[126][136]=0;
        ram[127][0]=0;ram[127][1]=1;ram[127][2]=0;ram[127][3]=1;ram[127][4]=0;ram[127][5]=1;ram[127][6]=1;ram[127][7]=1;ram[127][8]=0;ram[127][9]=1;ram[127][10]=1;ram[127][11]=1;ram[127][12]=1;ram[127][13]=1;ram[127][14]=1;ram[127][15]=1;ram[127][16]=1;ram[127][17]=1;ram[127][18]=1;ram[127][19]=0;ram[127][20]=0;ram[127][21]=1;ram[127][22]=0;ram[127][23]=1;ram[127][24]=1;ram[127][25]=0;ram[127][26]=1;ram[127][27]=1;ram[127][28]=0;ram[127][29]=1;ram[127][30]=0;ram[127][31]=0;ram[127][32]=0;ram[127][33]=1;ram[127][34]=1;ram[127][35]=0;ram[127][36]=1;ram[127][37]=1;ram[127][38]=0;ram[127][39]=1;ram[127][40]=1;ram[127][41]=0;ram[127][42]=1;ram[127][43]=1;ram[127][44]=1;ram[127][45]=1;ram[127][46]=1;ram[127][47]=0;ram[127][48]=0;ram[127][49]=1;ram[127][50]=1;ram[127][51]=1;ram[127][52]=0;ram[127][53]=1;ram[127][54]=1;ram[127][55]=1;ram[127][56]=1;ram[127][57]=1;ram[127][58]=1;ram[127][59]=1;ram[127][60]=1;ram[127][61]=1;ram[127][62]=0;ram[127][63]=1;ram[127][64]=0;ram[127][65]=0;ram[127][66]=1;ram[127][67]=1;ram[127][68]=0;ram[127][69]=1;ram[127][70]=0;ram[127][71]=0;ram[127][72]=1;ram[127][73]=1;ram[127][74]=1;ram[127][75]=1;ram[127][76]=1;ram[127][77]=1;ram[127][78]=0;ram[127][79]=0;ram[127][80]=1;ram[127][81]=1;ram[127][82]=0;ram[127][83]=1;ram[127][84]=0;ram[127][85]=0;ram[127][86]=0;ram[127][87]=0;ram[127][88]=1;ram[127][89]=1;ram[127][90]=1;ram[127][91]=1;ram[127][92]=0;ram[127][93]=1;ram[127][94]=0;ram[127][95]=0;ram[127][96]=1;ram[127][97]=1;ram[127][98]=1;ram[127][99]=1;ram[127][100]=1;ram[127][101]=0;ram[127][102]=0;ram[127][103]=1;ram[127][104]=1;ram[127][105]=1;ram[127][106]=0;ram[127][107]=1;ram[127][108]=1;ram[127][109]=1;ram[127][110]=1;ram[127][111]=1;ram[127][112]=1;ram[127][113]=0;ram[127][114]=1;ram[127][115]=0;ram[127][116]=0;ram[127][117]=1;ram[127][118]=1;ram[127][119]=1;ram[127][120]=0;ram[127][121]=1;ram[127][122]=1;ram[127][123]=0;ram[127][124]=0;ram[127][125]=1;ram[127][126]=0;ram[127][127]=1;ram[127][128]=0;ram[127][129]=0;ram[127][130]=1;ram[127][131]=1;ram[127][132]=1;ram[127][133]=0;ram[127][134]=0;ram[127][135]=1;ram[127][136]=1;
        ram[128][0]=0;ram[128][1]=1;ram[128][2]=1;ram[128][3]=1;ram[128][4]=1;ram[128][5]=0;ram[128][6]=1;ram[128][7]=0;ram[128][8]=1;ram[128][9]=1;ram[128][10]=0;ram[128][11]=0;ram[128][12]=1;ram[128][13]=1;ram[128][14]=1;ram[128][15]=0;ram[128][16]=1;ram[128][17]=1;ram[128][18]=1;ram[128][19]=1;ram[128][20]=1;ram[128][21]=1;ram[128][22]=1;ram[128][23]=1;ram[128][24]=1;ram[128][25]=0;ram[128][26]=1;ram[128][27]=0;ram[128][28]=1;ram[128][29]=1;ram[128][30]=1;ram[128][31]=1;ram[128][32]=0;ram[128][33]=1;ram[128][34]=0;ram[128][35]=1;ram[128][36]=0;ram[128][37]=1;ram[128][38]=1;ram[128][39]=0;ram[128][40]=1;ram[128][41]=0;ram[128][42]=0;ram[128][43]=0;ram[128][44]=0;ram[128][45]=0;ram[128][46]=0;ram[128][47]=0;ram[128][48]=0;ram[128][49]=1;ram[128][50]=0;ram[128][51]=1;ram[128][52]=1;ram[128][53]=0;ram[128][54]=0;ram[128][55]=0;ram[128][56]=1;ram[128][57]=1;ram[128][58]=1;ram[128][59]=1;ram[128][60]=0;ram[128][61]=1;ram[128][62]=0;ram[128][63]=0;ram[128][64]=0;ram[128][65]=1;ram[128][66]=1;ram[128][67]=1;ram[128][68]=1;ram[128][69]=0;ram[128][70]=0;ram[128][71]=1;ram[128][72]=0;ram[128][73]=1;ram[128][74]=0;ram[128][75]=0;ram[128][76]=1;ram[128][77]=0;ram[128][78]=1;ram[128][79]=1;ram[128][80]=1;ram[128][81]=1;ram[128][82]=1;ram[128][83]=1;ram[128][84]=1;ram[128][85]=1;ram[128][86]=0;ram[128][87]=1;ram[128][88]=1;ram[128][89]=1;ram[128][90]=1;ram[128][91]=0;ram[128][92]=1;ram[128][93]=1;ram[128][94]=1;ram[128][95]=1;ram[128][96]=0;ram[128][97]=1;ram[128][98]=0;ram[128][99]=1;ram[128][100]=1;ram[128][101]=1;ram[128][102]=1;ram[128][103]=0;ram[128][104]=1;ram[128][105]=0;ram[128][106]=1;ram[128][107]=0;ram[128][108]=1;ram[128][109]=1;ram[128][110]=0;ram[128][111]=0;ram[128][112]=0;ram[128][113]=1;ram[128][114]=1;ram[128][115]=0;ram[128][116]=1;ram[128][117]=1;ram[128][118]=0;ram[128][119]=0;ram[128][120]=0;ram[128][121]=0;ram[128][122]=1;ram[128][123]=1;ram[128][124]=1;ram[128][125]=1;ram[128][126]=0;ram[128][127]=1;ram[128][128]=1;ram[128][129]=0;ram[128][130]=0;ram[128][131]=0;ram[128][132]=1;ram[128][133]=0;ram[128][134]=0;ram[128][135]=1;ram[128][136]=0;
        ram[129][0]=1;ram[129][1]=0;ram[129][2]=0;ram[129][3]=1;ram[129][4]=1;ram[129][5]=1;ram[129][6]=0;ram[129][7]=0;ram[129][8]=1;ram[129][9]=1;ram[129][10]=0;ram[129][11]=0;ram[129][12]=1;ram[129][13]=1;ram[129][14]=1;ram[129][15]=1;ram[129][16]=0;ram[129][17]=1;ram[129][18]=1;ram[129][19]=1;ram[129][20]=0;ram[129][21]=0;ram[129][22]=0;ram[129][23]=1;ram[129][24]=1;ram[129][25]=0;ram[129][26]=1;ram[129][27]=1;ram[129][28]=0;ram[129][29]=1;ram[129][30]=1;ram[129][31]=1;ram[129][32]=0;ram[129][33]=1;ram[129][34]=0;ram[129][35]=0;ram[129][36]=1;ram[129][37]=1;ram[129][38]=1;ram[129][39]=1;ram[129][40]=1;ram[129][41]=1;ram[129][42]=0;ram[129][43]=0;ram[129][44]=0;ram[129][45]=1;ram[129][46]=1;ram[129][47]=1;ram[129][48]=1;ram[129][49]=1;ram[129][50]=0;ram[129][51]=1;ram[129][52]=0;ram[129][53]=0;ram[129][54]=1;ram[129][55]=1;ram[129][56]=1;ram[129][57]=1;ram[129][58]=0;ram[129][59]=1;ram[129][60]=1;ram[129][61]=1;ram[129][62]=1;ram[129][63]=0;ram[129][64]=1;ram[129][65]=1;ram[129][66]=1;ram[129][67]=0;ram[129][68]=1;ram[129][69]=1;ram[129][70]=1;ram[129][71]=1;ram[129][72]=1;ram[129][73]=0;ram[129][74]=0;ram[129][75]=1;ram[129][76]=1;ram[129][77]=1;ram[129][78]=1;ram[129][79]=0;ram[129][80]=1;ram[129][81]=1;ram[129][82]=1;ram[129][83]=1;ram[129][84]=1;ram[129][85]=0;ram[129][86]=1;ram[129][87]=1;ram[129][88]=1;ram[129][89]=0;ram[129][90]=0;ram[129][91]=1;ram[129][92]=1;ram[129][93]=0;ram[129][94]=0;ram[129][95]=0;ram[129][96]=0;ram[129][97]=1;ram[129][98]=1;ram[129][99]=1;ram[129][100]=1;ram[129][101]=0;ram[129][102]=1;ram[129][103]=1;ram[129][104]=0;ram[129][105]=1;ram[129][106]=1;ram[129][107]=1;ram[129][108]=1;ram[129][109]=1;ram[129][110]=1;ram[129][111]=1;ram[129][112]=0;ram[129][113]=0;ram[129][114]=1;ram[129][115]=1;ram[129][116]=0;ram[129][117]=1;ram[129][118]=1;ram[129][119]=1;ram[129][120]=0;ram[129][121]=1;ram[129][122]=1;ram[129][123]=0;ram[129][124]=0;ram[129][125]=0;ram[129][126]=0;ram[129][127]=1;ram[129][128]=0;ram[129][129]=0;ram[129][130]=0;ram[129][131]=1;ram[129][132]=1;ram[129][133]=1;ram[129][134]=1;ram[129][135]=1;ram[129][136]=0;
        ram[130][0]=0;ram[130][1]=1;ram[130][2]=0;ram[130][3]=0;ram[130][4]=1;ram[130][5]=1;ram[130][6]=0;ram[130][7]=1;ram[130][8]=0;ram[130][9]=0;ram[130][10]=1;ram[130][11]=0;ram[130][12]=1;ram[130][13]=1;ram[130][14]=1;ram[130][15]=0;ram[130][16]=1;ram[130][17]=0;ram[130][18]=0;ram[130][19]=0;ram[130][20]=1;ram[130][21]=1;ram[130][22]=1;ram[130][23]=1;ram[130][24]=1;ram[130][25]=1;ram[130][26]=0;ram[130][27]=1;ram[130][28]=1;ram[130][29]=1;ram[130][30]=0;ram[130][31]=1;ram[130][32]=1;ram[130][33]=1;ram[130][34]=1;ram[130][35]=0;ram[130][36]=1;ram[130][37]=0;ram[130][38]=1;ram[130][39]=0;ram[130][40]=0;ram[130][41]=1;ram[130][42]=1;ram[130][43]=1;ram[130][44]=1;ram[130][45]=1;ram[130][46]=1;ram[130][47]=1;ram[130][48]=1;ram[130][49]=0;ram[130][50]=0;ram[130][51]=1;ram[130][52]=0;ram[130][53]=1;ram[130][54]=1;ram[130][55]=0;ram[130][56]=1;ram[130][57]=1;ram[130][58]=0;ram[130][59]=1;ram[130][60]=0;ram[130][61]=1;ram[130][62]=1;ram[130][63]=0;ram[130][64]=0;ram[130][65]=0;ram[130][66]=0;ram[130][67]=1;ram[130][68]=1;ram[130][69]=1;ram[130][70]=1;ram[130][71]=1;ram[130][72]=1;ram[130][73]=1;ram[130][74]=0;ram[130][75]=1;ram[130][76]=1;ram[130][77]=1;ram[130][78]=0;ram[130][79]=0;ram[130][80]=1;ram[130][81]=0;ram[130][82]=1;ram[130][83]=0;ram[130][84]=1;ram[130][85]=1;ram[130][86]=1;ram[130][87]=1;ram[130][88]=1;ram[130][89]=1;ram[130][90]=1;ram[130][91]=1;ram[130][92]=0;ram[130][93]=0;ram[130][94]=1;ram[130][95]=1;ram[130][96]=1;ram[130][97]=0;ram[130][98]=1;ram[130][99]=1;ram[130][100]=1;ram[130][101]=1;ram[130][102]=0;ram[130][103]=0;ram[130][104]=1;ram[130][105]=1;ram[130][106]=1;ram[130][107]=1;ram[130][108]=1;ram[130][109]=1;ram[130][110]=0;ram[130][111]=1;ram[130][112]=1;ram[130][113]=1;ram[130][114]=1;ram[130][115]=0;ram[130][116]=0;ram[130][117]=1;ram[130][118]=0;ram[130][119]=0;ram[130][120]=1;ram[130][121]=1;ram[130][122]=1;ram[130][123]=0;ram[130][124]=1;ram[130][125]=0;ram[130][126]=0;ram[130][127]=1;ram[130][128]=1;ram[130][129]=1;ram[130][130]=0;ram[130][131]=0;ram[130][132]=0;ram[130][133]=1;ram[130][134]=0;ram[130][135]=0;ram[130][136]=1;
        ram[131][0]=1;ram[131][1]=1;ram[131][2]=0;ram[131][3]=1;ram[131][4]=0;ram[131][5]=0;ram[131][6]=1;ram[131][7]=1;ram[131][8]=1;ram[131][9]=1;ram[131][10]=0;ram[131][11]=1;ram[131][12]=1;ram[131][13]=1;ram[131][14]=0;ram[131][15]=0;ram[131][16]=1;ram[131][17]=1;ram[131][18]=1;ram[131][19]=0;ram[131][20]=1;ram[131][21]=1;ram[131][22]=1;ram[131][23]=0;ram[131][24]=0;ram[131][25]=1;ram[131][26]=0;ram[131][27]=1;ram[131][28]=1;ram[131][29]=1;ram[131][30]=1;ram[131][31]=1;ram[131][32]=0;ram[131][33]=0;ram[131][34]=0;ram[131][35]=1;ram[131][36]=1;ram[131][37]=1;ram[131][38]=1;ram[131][39]=1;ram[131][40]=1;ram[131][41]=1;ram[131][42]=0;ram[131][43]=0;ram[131][44]=0;ram[131][45]=1;ram[131][46]=1;ram[131][47]=1;ram[131][48]=1;ram[131][49]=1;ram[131][50]=1;ram[131][51]=1;ram[131][52]=0;ram[131][53]=0;ram[131][54]=0;ram[131][55]=0;ram[131][56]=0;ram[131][57]=1;ram[131][58]=1;ram[131][59]=0;ram[131][60]=1;ram[131][61]=1;ram[131][62]=1;ram[131][63]=0;ram[131][64]=1;ram[131][65]=1;ram[131][66]=1;ram[131][67]=0;ram[131][68]=1;ram[131][69]=0;ram[131][70]=1;ram[131][71]=1;ram[131][72]=0;ram[131][73]=1;ram[131][74]=1;ram[131][75]=0;ram[131][76]=1;ram[131][77]=0;ram[131][78]=1;ram[131][79]=1;ram[131][80]=1;ram[131][81]=1;ram[131][82]=1;ram[131][83]=1;ram[131][84]=1;ram[131][85]=0;ram[131][86]=1;ram[131][87]=1;ram[131][88]=1;ram[131][89]=1;ram[131][90]=1;ram[131][91]=1;ram[131][92]=0;ram[131][93]=1;ram[131][94]=1;ram[131][95]=0;ram[131][96]=1;ram[131][97]=1;ram[131][98]=0;ram[131][99]=1;ram[131][100]=0;ram[131][101]=1;ram[131][102]=1;ram[131][103]=0;ram[131][104]=0;ram[131][105]=1;ram[131][106]=0;ram[131][107]=1;ram[131][108]=1;ram[131][109]=1;ram[131][110]=1;ram[131][111]=0;ram[131][112]=1;ram[131][113]=0;ram[131][114]=1;ram[131][115]=0;ram[131][116]=1;ram[131][117]=1;ram[131][118]=1;ram[131][119]=1;ram[131][120]=1;ram[131][121]=1;ram[131][122]=1;ram[131][123]=0;ram[131][124]=1;ram[131][125]=1;ram[131][126]=1;ram[131][127]=1;ram[131][128]=1;ram[131][129]=0;ram[131][130]=0;ram[131][131]=1;ram[131][132]=0;ram[131][133]=0;ram[131][134]=0;ram[131][135]=1;ram[131][136]=1;
        ram[132][0]=1;ram[132][1]=1;ram[132][2]=0;ram[132][3]=0;ram[132][4]=0;ram[132][5]=1;ram[132][6]=0;ram[132][7]=0;ram[132][8]=1;ram[132][9]=0;ram[132][10]=0;ram[132][11]=0;ram[132][12]=0;ram[132][13]=1;ram[132][14]=0;ram[132][15]=1;ram[132][16]=1;ram[132][17]=0;ram[132][18]=1;ram[132][19]=1;ram[132][20]=0;ram[132][21]=1;ram[132][22]=1;ram[132][23]=1;ram[132][24]=1;ram[132][25]=1;ram[132][26]=1;ram[132][27]=1;ram[132][28]=1;ram[132][29]=0;ram[132][30]=0;ram[132][31]=0;ram[132][32]=1;ram[132][33]=1;ram[132][34]=1;ram[132][35]=1;ram[132][36]=1;ram[132][37]=0;ram[132][38]=1;ram[132][39]=1;ram[132][40]=1;ram[132][41]=0;ram[132][42]=1;ram[132][43]=0;ram[132][44]=1;ram[132][45]=1;ram[132][46]=1;ram[132][47]=1;ram[132][48]=0;ram[132][49]=1;ram[132][50]=0;ram[132][51]=0;ram[132][52]=1;ram[132][53]=0;ram[132][54]=0;ram[132][55]=1;ram[132][56]=1;ram[132][57]=1;ram[132][58]=1;ram[132][59]=1;ram[132][60]=0;ram[132][61]=1;ram[132][62]=0;ram[132][63]=0;ram[132][64]=0;ram[132][65]=1;ram[132][66]=1;ram[132][67]=1;ram[132][68]=0;ram[132][69]=0;ram[132][70]=0;ram[132][71]=0;ram[132][72]=1;ram[132][73]=1;ram[132][74]=1;ram[132][75]=1;ram[132][76]=1;ram[132][77]=1;ram[132][78]=1;ram[132][79]=1;ram[132][80]=1;ram[132][81]=0;ram[132][82]=0;ram[132][83]=1;ram[132][84]=1;ram[132][85]=1;ram[132][86]=0;ram[132][87]=1;ram[132][88]=0;ram[132][89]=0;ram[132][90]=1;ram[132][91]=1;ram[132][92]=1;ram[132][93]=1;ram[132][94]=1;ram[132][95]=1;ram[132][96]=1;ram[132][97]=1;ram[132][98]=1;ram[132][99]=1;ram[132][100]=1;ram[132][101]=1;ram[132][102]=1;ram[132][103]=1;ram[132][104]=0;ram[132][105]=0;ram[132][106]=1;ram[132][107]=1;ram[132][108]=1;ram[132][109]=0;ram[132][110]=1;ram[132][111]=1;ram[132][112]=1;ram[132][113]=0;ram[132][114]=1;ram[132][115]=1;ram[132][116]=1;ram[132][117]=1;ram[132][118]=1;ram[132][119]=0;ram[132][120]=1;ram[132][121]=1;ram[132][122]=0;ram[132][123]=0;ram[132][124]=0;ram[132][125]=0;ram[132][126]=1;ram[132][127]=0;ram[132][128]=1;ram[132][129]=0;ram[132][130]=1;ram[132][131]=1;ram[132][132]=1;ram[132][133]=1;ram[132][134]=1;ram[132][135]=1;ram[132][136]=1;
        ram[133][0]=0;ram[133][1]=1;ram[133][2]=0;ram[133][3]=1;ram[133][4]=1;ram[133][5]=1;ram[133][6]=0;ram[133][7]=0;ram[133][8]=1;ram[133][9]=1;ram[133][10]=1;ram[133][11]=0;ram[133][12]=0;ram[133][13]=1;ram[133][14]=1;ram[133][15]=1;ram[133][16]=1;ram[133][17]=0;ram[133][18]=0;ram[133][19]=1;ram[133][20]=1;ram[133][21]=1;ram[133][22]=1;ram[133][23]=1;ram[133][24]=1;ram[133][25]=0;ram[133][26]=1;ram[133][27]=1;ram[133][28]=0;ram[133][29]=1;ram[133][30]=1;ram[133][31]=1;ram[133][32]=1;ram[133][33]=0;ram[133][34]=1;ram[133][35]=0;ram[133][36]=1;ram[133][37]=1;ram[133][38]=1;ram[133][39]=1;ram[133][40]=1;ram[133][41]=1;ram[133][42]=0;ram[133][43]=1;ram[133][44]=1;ram[133][45]=1;ram[133][46]=0;ram[133][47]=1;ram[133][48]=1;ram[133][49]=1;ram[133][50]=1;ram[133][51]=1;ram[133][52]=0;ram[133][53]=1;ram[133][54]=0;ram[133][55]=1;ram[133][56]=1;ram[133][57]=0;ram[133][58]=1;ram[133][59]=1;ram[133][60]=0;ram[133][61]=1;ram[133][62]=1;ram[133][63]=1;ram[133][64]=1;ram[133][65]=0;ram[133][66]=1;ram[133][67]=1;ram[133][68]=1;ram[133][69]=1;ram[133][70]=0;ram[133][71]=1;ram[133][72]=0;ram[133][73]=1;ram[133][74]=1;ram[133][75]=1;ram[133][76]=1;ram[133][77]=1;ram[133][78]=1;ram[133][79]=1;ram[133][80]=1;ram[133][81]=1;ram[133][82]=0;ram[133][83]=0;ram[133][84]=0;ram[133][85]=0;ram[133][86]=1;ram[133][87]=0;ram[133][88]=0;ram[133][89]=1;ram[133][90]=1;ram[133][91]=0;ram[133][92]=0;ram[133][93]=1;ram[133][94]=1;ram[133][95]=1;ram[133][96]=1;ram[133][97]=0;ram[133][98]=0;ram[133][99]=0;ram[133][100]=1;ram[133][101]=1;ram[133][102]=0;ram[133][103]=0;ram[133][104]=1;ram[133][105]=0;ram[133][106]=1;ram[133][107]=1;ram[133][108]=1;ram[133][109]=1;ram[133][110]=1;ram[133][111]=0;ram[133][112]=1;ram[133][113]=1;ram[133][114]=1;ram[133][115]=0;ram[133][116]=0;ram[133][117]=1;ram[133][118]=1;ram[133][119]=1;ram[133][120]=1;ram[133][121]=1;ram[133][122]=1;ram[133][123]=1;ram[133][124]=1;ram[133][125]=1;ram[133][126]=1;ram[133][127]=1;ram[133][128]=0;ram[133][129]=0;ram[133][130]=1;ram[133][131]=1;ram[133][132]=1;ram[133][133]=0;ram[133][134]=0;ram[133][135]=1;ram[133][136]=0;
        ram[134][0]=1;ram[134][1]=1;ram[134][2]=1;ram[134][3]=1;ram[134][4]=0;ram[134][5]=1;ram[134][6]=0;ram[134][7]=0;ram[134][8]=0;ram[134][9]=1;ram[134][10]=1;ram[134][11]=0;ram[134][12]=1;ram[134][13]=0;ram[134][14]=1;ram[134][15]=0;ram[134][16]=1;ram[134][17]=0;ram[134][18]=0;ram[134][19]=1;ram[134][20]=1;ram[134][21]=0;ram[134][22]=1;ram[134][23]=1;ram[134][24]=1;ram[134][25]=1;ram[134][26]=1;ram[134][27]=1;ram[134][28]=0;ram[134][29]=1;ram[134][30]=0;ram[134][31]=0;ram[134][32]=1;ram[134][33]=1;ram[134][34]=1;ram[134][35]=1;ram[134][36]=1;ram[134][37]=0;ram[134][38]=1;ram[134][39]=0;ram[134][40]=0;ram[134][41]=0;ram[134][42]=0;ram[134][43]=1;ram[134][44]=1;ram[134][45]=1;ram[134][46]=1;ram[134][47]=1;ram[134][48]=1;ram[134][49]=1;ram[134][50]=1;ram[134][51]=0;ram[134][52]=1;ram[134][53]=1;ram[134][54]=1;ram[134][55]=1;ram[134][56]=0;ram[134][57]=1;ram[134][58]=0;ram[134][59]=1;ram[134][60]=1;ram[134][61]=0;ram[134][62]=1;ram[134][63]=1;ram[134][64]=1;ram[134][65]=1;ram[134][66]=0;ram[134][67]=1;ram[134][68]=1;ram[134][69]=0;ram[134][70]=1;ram[134][71]=0;ram[134][72]=1;ram[134][73]=1;ram[134][74]=1;ram[134][75]=1;ram[134][76]=1;ram[134][77]=1;ram[134][78]=0;ram[134][79]=1;ram[134][80]=1;ram[134][81]=1;ram[134][82]=1;ram[134][83]=1;ram[134][84]=1;ram[134][85]=1;ram[134][86]=0;ram[134][87]=0;ram[134][88]=1;ram[134][89]=0;ram[134][90]=1;ram[134][91]=1;ram[134][92]=1;ram[134][93]=1;ram[134][94]=0;ram[134][95]=1;ram[134][96]=1;ram[134][97]=0;ram[134][98]=0;ram[134][99]=1;ram[134][100]=1;ram[134][101]=0;ram[134][102]=1;ram[134][103]=1;ram[134][104]=0;ram[134][105]=0;ram[134][106]=1;ram[134][107]=1;ram[134][108]=0;ram[134][109]=0;ram[134][110]=0;ram[134][111]=1;ram[134][112]=1;ram[134][113]=1;ram[134][114]=0;ram[134][115]=1;ram[134][116]=1;ram[134][117]=1;ram[134][118]=0;ram[134][119]=1;ram[134][120]=0;ram[134][121]=1;ram[134][122]=0;ram[134][123]=0;ram[134][124]=1;ram[134][125]=0;ram[134][126]=1;ram[134][127]=1;ram[134][128]=1;ram[134][129]=0;ram[134][130]=1;ram[134][131]=1;ram[134][132]=1;ram[134][133]=1;ram[134][134]=1;ram[134][135]=0;ram[134][136]=1;
        ram[135][0]=0;ram[135][1]=1;ram[135][2]=1;ram[135][3]=0;ram[135][4]=1;ram[135][5]=1;ram[135][6]=0;ram[135][7]=1;ram[135][8]=1;ram[135][9]=1;ram[135][10]=1;ram[135][11]=1;ram[135][12]=0;ram[135][13]=0;ram[135][14]=1;ram[135][15]=1;ram[135][16]=0;ram[135][17]=1;ram[135][18]=1;ram[135][19]=1;ram[135][20]=1;ram[135][21]=0;ram[135][22]=1;ram[135][23]=0;ram[135][24]=1;ram[135][25]=1;ram[135][26]=1;ram[135][27]=1;ram[135][28]=0;ram[135][29]=1;ram[135][30]=1;ram[135][31]=1;ram[135][32]=1;ram[135][33]=0;ram[135][34]=1;ram[135][35]=1;ram[135][36]=0;ram[135][37]=1;ram[135][38]=1;ram[135][39]=0;ram[135][40]=1;ram[135][41]=1;ram[135][42]=1;ram[135][43]=1;ram[135][44]=1;ram[135][45]=0;ram[135][46]=0;ram[135][47]=0;ram[135][48]=1;ram[135][49]=1;ram[135][50]=1;ram[135][51]=0;ram[135][52]=0;ram[135][53]=0;ram[135][54]=1;ram[135][55]=1;ram[135][56]=0;ram[135][57]=1;ram[135][58]=0;ram[135][59]=0;ram[135][60]=1;ram[135][61]=1;ram[135][62]=1;ram[135][63]=0;ram[135][64]=1;ram[135][65]=1;ram[135][66]=1;ram[135][67]=1;ram[135][68]=1;ram[135][69]=1;ram[135][70]=1;ram[135][71]=1;ram[135][72]=1;ram[135][73]=1;ram[135][74]=0;ram[135][75]=1;ram[135][76]=1;ram[135][77]=0;ram[135][78]=0;ram[135][79]=1;ram[135][80]=1;ram[135][81]=0;ram[135][82]=1;ram[135][83]=1;ram[135][84]=1;ram[135][85]=1;ram[135][86]=1;ram[135][87]=0;ram[135][88]=0;ram[135][89]=0;ram[135][90]=1;ram[135][91]=0;ram[135][92]=0;ram[135][93]=0;ram[135][94]=1;ram[135][95]=1;ram[135][96]=1;ram[135][97]=1;ram[135][98]=1;ram[135][99]=1;ram[135][100]=1;ram[135][101]=0;ram[135][102]=0;ram[135][103]=0;ram[135][104]=0;ram[135][105]=1;ram[135][106]=1;ram[135][107]=1;ram[135][108]=0;ram[135][109]=1;ram[135][110]=1;ram[135][111]=0;ram[135][112]=0;ram[135][113]=1;ram[135][114]=1;ram[135][115]=1;ram[135][116]=1;ram[135][117]=0;ram[135][118]=0;ram[135][119]=1;ram[135][120]=0;ram[135][121]=0;ram[135][122]=1;ram[135][123]=0;ram[135][124]=0;ram[135][125]=1;ram[135][126]=1;ram[135][127]=1;ram[135][128]=0;ram[135][129]=1;ram[135][130]=1;ram[135][131]=0;ram[135][132]=1;ram[135][133]=1;ram[135][134]=1;ram[135][135]=0;ram[135][136]=0;
        ram[136][0]=1;ram[136][1]=1;ram[136][2]=0;ram[136][3]=0;ram[136][4]=0;ram[136][5]=0;ram[136][6]=0;ram[136][7]=0;ram[136][8]=0;ram[136][9]=0;ram[136][10]=1;ram[136][11]=0;ram[136][12]=1;ram[136][13]=1;ram[136][14]=1;ram[136][15]=1;ram[136][16]=0;ram[136][17]=1;ram[136][18]=1;ram[136][19]=0;ram[136][20]=0;ram[136][21]=0;ram[136][22]=1;ram[136][23]=1;ram[136][24]=0;ram[136][25]=0;ram[136][26]=0;ram[136][27]=0;ram[136][28]=1;ram[136][29]=1;ram[136][30]=1;ram[136][31]=0;ram[136][32]=0;ram[136][33]=0;ram[136][34]=1;ram[136][35]=0;ram[136][36]=1;ram[136][37]=0;ram[136][38]=1;ram[136][39]=0;ram[136][40]=0;ram[136][41]=1;ram[136][42]=1;ram[136][43]=1;ram[136][44]=0;ram[136][45]=0;ram[136][46]=1;ram[136][47]=1;ram[136][48]=0;ram[136][49]=1;ram[136][50]=1;ram[136][51]=1;ram[136][52]=0;ram[136][53]=1;ram[136][54]=1;ram[136][55]=0;ram[136][56]=0;ram[136][57]=1;ram[136][58]=0;ram[136][59]=0;ram[136][60]=1;ram[136][61]=1;ram[136][62]=1;ram[136][63]=1;ram[136][64]=1;ram[136][65]=0;ram[136][66]=1;ram[136][67]=1;ram[136][68]=0;ram[136][69]=1;ram[136][70]=1;ram[136][71]=0;ram[136][72]=0;ram[136][73]=0;ram[136][74]=0;ram[136][75]=1;ram[136][76]=0;ram[136][77]=1;ram[136][78]=0;ram[136][79]=0;ram[136][80]=0;ram[136][81]=0;ram[136][82]=1;ram[136][83]=1;ram[136][84]=1;ram[136][85]=0;ram[136][86]=1;ram[136][87]=1;ram[136][88]=1;ram[136][89]=1;ram[136][90]=0;ram[136][91]=0;ram[136][92]=1;ram[136][93]=1;ram[136][94]=1;ram[136][95]=0;ram[136][96]=1;ram[136][97]=1;ram[136][98]=1;ram[136][99]=1;ram[136][100]=1;ram[136][101]=0;ram[136][102]=0;ram[136][103]=0;ram[136][104]=1;ram[136][105]=1;ram[136][106]=1;ram[136][107]=1;ram[136][108]=1;ram[136][109]=1;ram[136][110]=1;ram[136][111]=0;ram[136][112]=1;ram[136][113]=1;ram[136][114]=1;ram[136][115]=1;ram[136][116]=1;ram[136][117]=1;ram[136][118]=1;ram[136][119]=1;ram[136][120]=1;ram[136][121]=1;ram[136][122]=1;ram[136][123]=0;ram[136][124]=0;ram[136][125]=0;ram[136][126]=1;ram[136][127]=1;ram[136][128]=1;ram[136][129]=1;ram[136][130]=0;ram[136][131]=1;ram[136][132]=0;ram[136][133]=0;ram[136][134]=1;ram[136][135]=1;ram[136][136]=0;

        sum<=0;
    end
    
    genvar i;
    genvar j;
    generate
        for(i=0;i<size;i=i+1)
        begin: row
            for(j=0;j<size;j=j+1)
            begin: column
            
                if( (i==0 && (j==0 || j==size-1)) || (i==size-1 && (j==0 || j==size-1)) )
                begin: i_j_zero
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else sumram[i][j]=1;
                    end
                end
                
                else if(i==0)
                begin: i_zero
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else if (ram[i][j-1]+ram[i][j+1]+ram[i+1][j-1]+ram[i+1][j]+ram[i+1][j+1]<4)sumram[i][j]=1;
                        else sumram[i][j]=0;
                    end
                end
                
                else if(i==size-1)
                begin: i_end
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else if (ram[i][j-1]+ram[i][j+1]+ram[i-1][j-1]+ram[i-1][j]+ram[i-1][j+1]<4)sumram[i][j]=1;
                        else sumram[i][j]=0;
                    end
                end
                
                else if(j==0)
                begin: j_zero
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else if (ram[i-1][j]+ram[i-1][j+1]+ram[i][j+1]+ram[i+1][j]+ram[i+1][j+1]<4)sumram[i][j]=1;
                        else sumram[i][j]=0;
                    end
                end
                
                else if(j==size-1)
                begin: j_end
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else if (ram[i-1][j-1]+ram[i-1][j]+ram[i][j-1]+ram[i+1][j-1]+ram[i+1][j]<4)sumram[i][j]=1;
                        else sumram[i][j]=0;
                    end
                end
                
                else
                begin: normal
                    always @(*)
                    begin
                        if(rst||!ram[i][j])sumram[i][j]=0;
                        else if (ram[i-1][j-1]+ram[i-1][j]+ram[i-1][j+1]+ram[i][j-1]+ram[i][j+1]+ram[i+1][j-1]+ram[i+1][j]+ram[i+1][j+1]<4)sumram[i][j]=1;
                        else sumram[i][j]=0;
                    end
                end
            end
        end
    endgenerate
    
    integer c=0,d=0;
    reg [31:0]sum_cache=0;
    always @(*)
    begin
        sum_cache=0;
        for (c=0;c<size;c=c+1)
        begin: add_sumc
            for (d=0;d<size;d=d+1)
            begin: add_sumd
                sum_cache=sum_cache+sumram[c][d];
            end
        end
    end
        
    genvar a,b;
    generate
        for (a=0;a<size;a=a+1)
        begin: ram_row
            for (b=0;b<size;b=b+1)
            begin: ram_column
                always @(posedge clk) ram[a][b]<=ram[a][b]-sumram[a][b];
            end    
        end
    endgenerate
    
    always @(posedge clk)
    begin
        if(rst)sum<=0;
        else sum<=sum+sum_cache;
    end
    
endmodule

