`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09.01.2026 09:28:32
// Design Name: 
// Module Name: Main2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Main2(
    input clk,rst,
    output reg [63:0]ans
    );
    
    parameter size=194;
    
    reg [63:0]ram[2*size-1:0];
    initial
    begin
        ram[0]=64'd512859921084892;ram[1]=64'd514321322528165;ram[2]=64'd11256263100164;ram[3]=64'd12830604534729;ram[4]=64'd85116519420599;ram[5]=64'd87459851977631;ram[6]=64'd406717661663760;ram[7]=64'd407318544520029;ram[8]=64'd163452173268505;ram[9]=64'd163452173268505;ram[10]=64'd352163676002057;ram[11]=64'd353682906584490;ram[12]=64'd493917957460777;ram[13]=64'd499926818635595;ram[14]=64'd475214413811256;ram[15]=64'd475460418793114;ram[16]=64'd327589455877896;ram[17]=64'd330833236397342;ram[18]=64'd432793196663974;ram[19]=64'd438939090134058;ram[20]=64'd142021536452283;ram[21]=64'd142458197886533;ram[22]=64'd480576606153933;ram[23]=64'd481201233296425;ram[24]=64'd403027733769497;ram[25]=64'd403528723415276;ram[26]=64'd280425795751218;ram[27]=64'd280425795751218;ram[28]=64'd475543316179274;ram[29]=64'd475865041061127;ram[30]=64'd365311178187035;
        ram[31]=64'd371696619383403;ram[32]=64'd345195747812243;ram[33]=64'd348539598024039;ram[34]=64'd244367967651559;ram[35]=64'd246443094684012;ram[36]=64'd282225709715432;ram[37]=64'd288948158549589;ram[38]=64'd2866510385568;ram[39]=64'd8245528252945;ram[40]=64'd102842075080213;ram[41]=64'd103099712594499;ram[42]=64'd477891742632187;ram[43]=64'd478557346319753;ram[44]=64'd314471537564046;ram[45]=64'd318839025331372;ram[46]=64'd438939090134059;ram[47]=64'd438939090134059;ram[48]=64'd475543316179274;ram[49]=64'd475865041061127;ram[50]=64'd247597610136719;ram[51]=64'd249350770074688;ram[52]=64'd402391070936536;ram[53]=64'd403027733769497;ram[54]=64'd517440331784466;ram[55]=64'd518721200423551;ram[56]=64'd151853435379858;ram[57]=64'd159065340219307;ram[58]=64'd41365168848672;ram[59]=64'd41365168848672;ram[60]=64'd473192720395488;
        ram[61]=64'd473638033595403;ram[62]=64'd423459461472407;ram[63]=64'd428100785796806;ram[64]=64'd345195747812243;ram[65]=64'd348539598024039;ram[66]=64'd184720620231963;ram[67]=64'd189425282918814;ram[68]=64'd13437510189376;ram[69]=64'd14964953082632;ram[70]=64'd213043812181954;ram[71]=64'd216479274574897;ram[72]=64'd74729109838980;ram[73]=64'd79200808617434;ram[74]=64'd272402315102244;ram[75]=64'd280425795751218;ram[76]=64'd463372984834827;ram[77]=64'd469143037229218;ram[78]=64'd253435371892878;ram[79]=64'd259698393140249;ram[80]=64'd463372984834827;ram[81]=64'd469143037229218;ram[82]=64'd534250792816163;ram[83]=64'd541114169199412;ram[84]=64'd248846253931401;ram[85]=64'd250671481074223;ram[86]=64'd106618450507051;ram[87]=64'd107537813186427;ram[88]=64'd425223261695362;ram[89]=64'd430815552180428;ram[90]=64'd144221722700109;
        ram[91]=64'd144403316706296;ram[92]=64'd149447865448566;ram[93]=64'd149591163712297;ram[94]=64'd107537813186427;ram[95]=64'd108004960050726;ram[96]=64'd74729109838979;ram[97]=64'd74729109838979;ram[98]=64'd498638157843121;ram[99]=64'd499926818635595;ram[100]=64'd377723593244025;ram[101]=64'd381453006636276;ram[102]=64'd24469822545597;ram[103]=64'd28905036834526;ram[104]=64'd478959415634099;ram[105]=64'd479572266127678;ram[106]=64'd196631611793187;ram[107]=64'd199442731572520;ram[108]=64'd102601416161455;ram[109]=64'd103392608501004;ram[110]=64'd204293845440549;ram[111]=64'd204293845440549;ram[112]=64'd141942632584343;ram[113]=64'd142458197886533;ram[114]=64'd144403316706296;ram[115]=64'd144958336655671;ram[116]=64'd360271538394352;ram[117]=64'd361638424717532;ram[118]=64'd124327235911656;ram[119]=64'd128652000240528;ram[120]=64'd322478956945714;
        ram[121]=64'd330833236397342;ram[122]=64'd173143830650714;ram[123]=64'd177164492234604;ram[124]=64'd141548266176759;ram[125]=64'd141942632584343;ram[126]=64'd480182573513490;ram[127]=64'd480330678306927;ram[128]=64'd473760735647262;ram[129]=64'd474406582226503;ram[130]=64'd405329367317474;ram[131]=64'd406051406189253;ram[132]=64'd504270134722688;ram[133]=64'd512029242808107;ram[134]=64'd479475085586324;ram[135]=64'd479572266127678;ram[136]=64'd18426346679546;ram[137]=64'd19777543329085;ram[138]=64'd2866510385568;ram[139]=64'd4231745022169;ram[140]=64'd149591163712297;ram[141]=64'd149919936790602;ram[142]=64'd525604737586813;ram[143]=64'd528523145466224;ram[144]=64'd358987141008867;ram[145]=64'd360624439822697;ram[146]=64'd382516644929553;ram[147]=64'd388406164141792;ram[148]=64'd145331203961556;ram[149]=64'd146046820232156;ram[150]=64'd14237415584385;
        ram[151]=64'd15924049948423;ram[152]=64'd374209474121225;ram[153]=64'd377723593244023;ram[154]=64'd334687610529456;ram[155]=64'd335663735053582;ram[156]=64'd155033974759271;ram[157]=64'd157349828556626;ram[158]=64'd114366847962685;ram[159]=64'd116294965915693;ram[160]=64'd355930697101159;ram[161]=64'd357557290228042;ram[162]=64'd163452173268505;ram[163]=64'd170189020588494;ram[164]=64'd10200758506934;ram[165]=64'd11675873319750;ram[166]=64'd479882960182177;ram[167]=64'd480330678306927;ram[168]=64'd445042671814231;ram[169]=64'd445042671814231;ram[170]=64'd480330678306927;ram[171]=64'd480974894454623;ram[172]=64'd306258271480626;ram[173]=64'd307968155504989;ram[174]=64'd519398465210473;ram[175]=64'd520540738946159;ram[176]=64'd223229557785366;ram[177]=64'd227025154757080;ram[178]=64'd99488387218746;ram[179]=64'd99488387218746;ram[180]=64'd354062340382732;
        ram[181]=64'd355800257907019;ram[182]=64'd335663735053583;ram[183]=64'd339871336806922;ram[184]=64'd474035001338741;ram[185]=64'd474922781605310;ram[186]=64'd545078918614008;ram[187]=64'd547008360559588;ram[188]=64'd22317984096899;ram[189]=64'd26888145536722;ram[190]=64'd407085583465386;ram[191]=64'd407318544520029;ram[192]=64'd405568050903009;ram[193]=64'd406288084821195;ram[194]=64'd232046628549385;ram[195]=64'd239886267027114;ram[196]=64'd103392608501004;ram[197]=64'd104133217219567;ram[198]=64'd146046820232156;ram[199]=64'd146322411858073;ram[200]=64'd392975504911599;ram[201]=64'd400490540710331;ram[202]=64'd353016434053625;ram[203]=64'd354748246306487;ram[204]=64'd455335377063119;ram[205]=64'd457899212781249;ram[206]=64'd215156606188916;ram[207]=64'd219455334407782;ram[208]=64'd144403316706296;ram[209]=64'd145205574339865;ram[210]=64'd282225709715432;
        ram[211]=64'd286354786062902;ram[212]=64'd102493040223700;ram[213]=64'd102601416161455;ram[214]=64'd402654937231438;ram[215]=64'd403027733769497;ram[216]=64'd475460418793114;ram[217]=64'd476059605944812;ram[218]=64'd122091435294890;ram[219]=64'd124327235911654;ram[220]=64'd547008360559589;ram[221]=64'd552361753325632;ram[222]=64'd516690820098898;ram[223]=64'd517792845762147;ram[224]=64'd102601416161455;ram[225]=64'd103392608501004;ram[226]=64'd515515480200760;ram[227]=64'd517024089221025;ram[228]=64'd227025154757081;ram[229]=64'd228788136841922;ram[230]=64'd388406164141793;ram[231]=64'd388406164141793;ram[232]=64'd245731070582959;ram[233]=64'd247896713915077;ram[234]=64'd147682702289292;ram[235]=64'd147944111104358;ram[236]=64'd232046628549385;ram[237]=64'd236269038299131;ram[238]=64'd101727995252076;ram[239]=64'd101893597192742;ram[240]=64'd146322411858073;
        ram[241]=64'd146827505938482;ram[242]=64'd265768889540204;ram[243]=64'd268076557887533;ram[244]=64'd362644837883327;ram[245]=64'd369172553644526;ram[246]=64'd453347800747762;ram[247]=64'd460712954322341;ram[248]=64'd302023237296177;ram[249]=64'd311369101986143;ram[250]=64'd92074568264509;ram[251]=64'd99488387218745;ram[252]=64'd534250792816163;ram[253]=64'd538759869162311;ram[254]=64'd514644567422522;ram[255]=64'd516286219051199;ram[256]=64'd142021536452283;ram[257]=64'd142458197886533;ram[258]=64'd103099712594499;ram[259]=64'd103994931941778;ram[260]=64'd108661255859598;ram[261]=64'd108966250607200;ram[262]=64'd476782263335539;ram[263]=64'd477219301791520;ram[264]=64'd406288084821195;ram[265]=64'd406717661663760;ram[266]=64'd293049127369610;ram[267]=64'd300062402676600;ram[268]=64'd354947816816014;ram[269]=64'd356630527176192;ram[270]=64'd513863705373574;
        ram[271]=64'd515076772891135;ram[272]=64'd402654937231438;ram[273]=64'd403307611288314;ram[274]=64'd35269914317143;ram[275]=64'd39695782939342;ram[276]=64'd148889419672007;ram[277]=64'd149591163712297;ram[278]=64'd242798507145598;ram[279]=64'd245493573576481;ram[280]=64'd520076800433250;ram[281]=64'd521519731841702;ram[282]=64'd105125698669905;ram[283]=64'd105636844019680;ram[284]=64'd149919936790602;ram[285]=64'd150462928965633;ram[286]=64'd445042671814231;ram[287]=64'd451161917293972;ram[288]=64'd475214413811256;ram[289]=64'd475865041061127;ram[290]=64'd15184860973332;ram[291]=64'd16841529948392;ram[292]=64'd241575901323241;ram[293]=64'd243667417822264;ram[294]=64'd116294965915693;ram[295]=64'd116294965915693;ram[296]=64'd142021536452283;ram[297]=64'd142696958243488;ram[298]=64'd409976406315634;ram[299]=64'd410555272379186;ram[300]=64'd109214419527261;
        ram[301]=64'd109599415788054;ram[302]=64'd486282179063049;ram[303]=64'd491061824835978;ram[304]=64'd103099712594499;ram[305]=64'd103723767650008;ram[306]=64'd293049127369610;ram[307]=64'd293049127369610;ram[308]=64'd62226970078581;ram[309]=64'd69495982987098;ram[310]=64'd146322411858073;ram[311]=64'd146827505938482;ram[312]=64'd491061824835978;ram[313]=64'd491061824835978;ram[314]=64'd17179233651851;ram[315]=64'd18830111267124;ram[316]=64'd102493040223700;ram[317]=64'd102601416161455;ram[318]=64'd193866729256721;ram[319]=64'd199442731572520;ram[320]=64'd150212077211861;ram[321]=64'd150462928965633;ram[322]=64'd62226970078581;ram[323]=64'd69495982987098;ram[324]=64'd555240684135726;ram[325]=64'd560251920336867;ram[326]=64'd392975504911598;ram[327]=64'd392975504911598;ram[328]=64'd103723767650008;ram[329]=64'd104402500724508;ram[330]=64'd53992525017805;
        ram[331]=64'd58576571790780;ram[332]=64'd173143830650714;ram[333]=64'd177164492234604;ram[334]=64'd358291972543663;ram[335]=64'd359472466194581;ram[336]=64'd101228998017649;ram[337]=64'd101430434873838;ram[338]=64'd31655863277653;ram[339]=64'd35269914317142;ram[340]=64'd410315459676065;ram[341]=64'd410555272379186;ram[342]=64'd418544898567771;ram[343]=64'd418544898567771;ram[344]=64'd357209901292816;ram[345]=64'd358824045906136;ram[346]=64'd259698393140250;ram[347]=64'd259698393140250;ram[348]=64'd100960550591037;ram[349]=64'd101430434873838;ram[350]=64'd105636844019680;ram[351]=64'd106516704612369;ram[352]=64'd12449698691637;ram[353]=64'd13694195772711;ram[354]=64'd478387779303792;ram[355]=64'd479096686553970;ram[356]=64'd132729578205911;ram[357]=64'd136390389715745;ram[358]=64'd41365168848672;ram[359]=64'd49031435034747;ram[360]=64'd182050206515811;
        ram[361]=64'd184720620231961;ram[362]=64'd80798010743456;ram[363]=64'd89758941577635;ram[364]=64'd555240684135725;ram[365]=64'd555240684135725;ram[366]=64'd477219301791520;ram[367]=64'd477451665942660;ram[368]=64'd16284281899664;ram[369]=64'd18043423892091;ram[370]=64'd521077678197487;ram[371]=64'd522434838851811;ram[372]=64'd528523145466226;ram[373]=64'd529811726976053;ram[374]=64'd478092010393383;ram[375]=64'd478557346319753;ram[376]=64'd518551031596939;ram[377]=64'd519651768836269;ram[378]=64'd51716793013563;ram[379]=64'd58576571790780;ram[380]=64'd416293147622133;ram[381]=64'd418544898567771;ram[382]=64'd204293845440550;ram[383]=64'd209480228080573;ram[384]=64'd475865041061127;ram[385]=64'd476366294808733;ram[386]=64'd142458197886533;ram[387]=64'd142780858100993;
        ans=0;
    end
    
    //Sorting
    reg sort_decide=0; 
    always @(posedge clk) sort_decide<=~sort_decide;
    
    reg [31:0]j=0;
    reg [31:0]k=0;
    reg change=0;
    reg [31:0]start=0;
    reg [2:0]state=0;

    genvar i;
    generate
        for(i=0;i<2*size;i=i+2)
        begin: sorter
            always @(posedge clk)
            begin
                if(j==i && change)ram[i+1]<=ram[k+1];
                if(i%4)
                begin
                    if (sort_decide)
                    begin
                        if (ram[i]<ram[i-2])
                        begin
                            ram[i]<=ram[i-2];
                            ram[i+1]<=ram[i-1];
                        end
                        else if (ram[i]==ram[i-2] && ram[i-1]<ram[i+1])
                            ram[i+1]<=ram[i-1];
                    end
                    else
                    begin
                        if(i<2*size-2)
                        begin
                            if (ram[i]>ram[i+2])
                            begin
                                ram[i]<=ram[i+2];
                                ram[i+1]<=ram[i+3];
                            end
                            else if (ram[i]==ram[i+2] && ram[i+1]<ram[i+3])
                                ram[i+1]<=ram[i+3];
                        end
                    end
                end
                else
                begin
                    if (sort_decide)
                    begin
                        if (ram[i]>ram[i+2])
                        begin
                            ram[i]<=ram[i+2];
                            ram[i+1]<=ram[i+3];
                        end
                        else if (ram[i]==ram[i+2] && ram[i+1]<ram[i+3])
                            ram[i+1]<=ram[i+3];
                    end
                    else
                    begin
                        if(i<2*size-2)
                        begin
                            if (ram[i]<ram[i-2])
                            begin
                                ram[i]<=ram[i-2];
                                ram[i+1]<=ram[i-1];
                            end
                            else if (ram[i]==ram[i-2] && ram[i+1]>ram[i-1])
                                ram[i+1]<=ram[i-1];
                        end
                    end
                end
            end
        end
    endgenerate
    
    reg [63:0]max=0;
    always @(posedge clk)
    begin
        if(rst)
        begin
            j<=0;k<=0;start<=0;state<=0;change<=0;
            max<=ram[0];ans<=0;
        end
        else
        begin
            case(state)
            0:begin
                if(start<size)start<=start+1;
                else state<=1;
            end
            1:begin
                if(change)change<=0;
                else
                begin
                    if(k<2*size-2)
                    begin
                        k<=k+2;
                        if (ram[j]!=ram[k+2])
                        begin
                            if (ram[k+2]>ram[j+1]) j<=j+2;
                            else if (ram[j+1]<ram[k+3])change<=1;    
                        end
                    end   
                    else 
                    begin
                        state<=2;
                        k<=0;
                    end
                end
            end
            2:
            begin
                if(k<2*size)
                begin
                    k<=k+1;
                    if (!k[0] && ram[k]>=max)max<=ram[k];
                    else if (ram[k]>=max)
                    begin
                        ans<=ans+ram[k]-max+1;
                        max<=ram[k]+1;
                    end
                end
            end
            endcase
        end
    end
endmodule
