`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.01.2026 22:31:24
// Design Name: 
// Module Name: Main1_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Main1_tb();
    reg clk,rst;
    reg [63:0]ip;
    wire [15:0]ans;
    
    Main1 DUT(
        .clk(clk),
        .rst(rst),
        .ip(ip),
        .ans(ans)
    );

    always #5 clk=~clk;
    
    initial
    begin
        clk=0;rst=0;ip=0;
        #10;
        ip=64'd329928111646776;#10;ip=64'd482309026155231;#10;ip=64'd525241827868042;#10;ip=64'd96135717389080;#10;ip=64'd499110589511466;#10;ip=64'd308522093992965;#10;ip=64'd33674948675734;#10;ip=64'd430565826580167;#10;ip=64'd414408953001629;#10;ip=64'd173680629421068;#10;ip=64'd548677463098858;#10;ip=64'd494697327482911;#10;ip=64'd206935857962233;#10;ip=64'd288752505984903;#10;ip=64'd316429280970249;#10;ip=64'd495713402865828;#10;ip=64'd169490817148712;#10;ip=64'd368483521093476;#10;ip=64'd258261134664607;#10;ip=64'd495149959285654;#10;ip=64'd475606183862234;#10;ip=64'd305251526450866;#10;ip=64'd225901258916804;#10;ip=64'd445966182017246;#10;ip=64'd434250874173072;#10;ip=64'd82915457820367;#10;ip=64'd97393274258734;#10;ip=64'd285494998420898;#10;ip=64'd502528740343165;#10;ip=64'd274566425378261;#10;ip=64'd470846785856273;#10;ip=64'd136708479249460;#10;ip=64'd162283218276275;#10;ip=64'd393591452022683;#10;ip=64'd460376379554779;#10;ip=64'd105696714402057;#10;ip=64'd511104696139372;#10;ip=64'd351529171768347;#10;ip=64'd547381378685144;#10;ip=64'd68431490253071;#10;ip=64'd298153102009441;#10;ip=64'd85916336633004;#10;ip=64'd66955289166933;#10;ip=64'd407098341285956;#10;ip=64'd542255776457073;#10;ip=64'd508930162141684;#10;ip=64'd66827379778215;#10;ip=64'd279783855088048;#10;ip=64'd492398265075615;#10;ip=64'd248767410738826;#10;ip=64'd197872398759823;#10;ip=64'd143340810943871;#10;ip=64'd46011637170446;#10;ip=64'd126524553899277;#10;ip=64'd156815771597592;#10;ip=64'd452835811023038;#10;ip=64'd274204463983422;#10;ip=64'd255067341756469;#10;ip=64'd540234469303121;#10;ip=64'd496987139396868;#10;ip=64'd555891985373714;#10;ip=64'd225388263513271;#10;ip=64'd262459661861113;#10;ip=64'd87225975280979;#10;ip=64'd53720559983785;#10;ip=64'd177882066763557;#10;ip=64'd288801648898790;#10;ip=64'd63791472295914;#10;ip=64'd352250011831260;#10;ip=64'd206278464247171;#10;ip=64'd134788841536024;#10;ip=64'd335032464310109;#10;ip=64'd556514653083429;#10;ip=64'd413516863406264;#10;ip=64'd161347101973576;#10;ip=64'd545399029770191;#10;ip=64'd472829659788930;#10;ip=64'd360231799823876;#10;ip=64'd156760218821562;#10;ip=64'd75012555232544;#10;ip=64'd189163976519132;#10;ip=64'd305431230444124;#10;ip=64'd47556076381637;#10;ip=64'd484236835622830;#10;ip=64'd323037782466288;#10;ip=64'd248260546770241;#10;ip=64'd385916685909473;#10;ip=64'd176553924738469;#10;ip=64'd315979862702759;#10;ip=64'd427290550436004;#10;ip=64'd437046249326037;#10;ip=64'd107897638650226;#10;ip=64'd173287681178617;#10;ip=64'd377567155948386;#10;ip=64'd23821440169790;#10;ip=64'd455789236975611;#10;ip=64'd468616497372607;#10;ip=64'd351630682027145;#10;ip=64'd475247397314142;#10;ip=64'd296694806740658;#10;ip=64'd400260298743488;#10;
        ip=64'd117829241442811;#10;ip=64'd530564276123775;#10;ip=64'd410991765233531;#10;ip=64'd462937925726291;#10;ip=64'd538975155010245;#10;ip=64'd94811163103973;#10;ip=64'd213777020819769;#10;ip=64'd266124223822590;#10;ip=64'd382897409024790;#10;ip=64'd389684560259599;#10;ip=64'd520301184003705;#10;ip=64'd14159977777584;#10;ip=64'd104526729594809;#10;ip=64'd265414483809986;#10;ip=64'd305160027113765;#10;ip=64'd145137875095728;#10;ip=64'd314789183106976;#10;ip=64'd84671645010572;#10;ip=64'd551192788962037;#10;ip=64'd63140952781035;#10;ip=64'd152790791169992;#10;ip=64'd358249314650523;#10;ip=64'd57619396015514;#10;ip=64'd371048477263502;#10;ip=64'd43723010091329;#10;ip=64'd354833015197434;#10;ip=64'd528978055728588;#10;ip=64'd397085006618713;#10;ip=64'd213967361863856;#10;ip=64'd359981491037828;#10;ip=64'd385991394542590;#10;ip=64'd259384895073422;#10;ip=64'd305382934938356;#10;ip=64'd325799054815220;#10;ip=64'd338355547018775;#10;ip=64'd385559913028576;#10;ip=64'd2197336567346;#10;ip=64'd186417713031811;#10;ip=64'd139160151867234;#10;ip=64'd345213498738360;#10;ip=64'd148218489601903;#10;ip=64'd371588279621791;#10;ip=64'd338635552506598;#10;ip=64'd96354674957257;#10;ip=64'd457655392901609;#10;ip=64'd68051467604790;#10;ip=64'd245777062929041;#10;ip=64'd93057662802800;#10;ip=64'd313438892416489;#10;ip=64'd417740659571195;#10;ip=64'd529072878715424;#10;ip=64'd120134767192617;#10;ip=64'd412091961105487;#10;ip=64'd106935868378177;#10;ip=64'd522069743249636;#10;ip=64'd260388524020154;#10;ip=64'd111666973903629;#10;ip=64'd44268407405977;#10;ip=64'd115572039812179;#10;ip=64'd293867232815220;#10;ip=64'd237260942030335;#10;ip=64'd246627332244583;#10;ip=64'd458113909274192;#10;ip=64'd557550691169619;#10;ip=64'd360390031192940;#10;ip=64'd166068283210014;#10;ip=64'd40963467930318;#10;ip=64'd342656301747653;#10;ip=64'd484652751523921;#10;ip=64'd92914650194336;#10;ip=64'd552705707274281;#10;ip=64'd193219271862351;#10;ip=64'd224135805639407;#10;ip=64'd450506060399134;#10;ip=64'd440031713484081;#10;ip=64'd296624565350139;#10;ip=64'd285148757973257;#10;ip=64'd317571583672140;#10;ip=64'd554270807901887;#10;ip=64'd427545994287941;#10;ip=64'd467886679084771;#10;ip=64'd20467538103182;#10;ip=64'd258043783652238;#10;ip=64'd31979007483159;#10;ip=64'd53914464635930;#10;ip=64'd67291764735355;#10;ip=64'd548056993839685;#10;ip=64'd145940474692981;#10;ip=64'd492618818691046;#10;ip=64'd543898596804083;#10;ip=64'd285079558926647;#10;ip=64'd266939889945458;#10;ip=64'd319144605258498;#10;ip=64'd82161508442190;#10;ip=64'd304656547859574;#10;ip=64'd333243314874982;#10;ip=64'd76620959106542;#10;ip=64'd447041570162937;#10;ip=64'd458031244195180;#10;ip=64'd196007380612049;#10;
        ip=64'd188668742770737;#10;ip=64'd301677694030334;#10;ip=64'd119718025553867;#10;ip=64'd65434272539891;#10;ip=64'd526378244569942;#10;ip=64'd299379972173118;#10;ip=64'd547393330166250;#10;ip=64'd149497804485190;#10;ip=64'd30730425184500;#10;ip=64'd125490524594151;#10;ip=64'd25511461942913;#10;ip=64'd542579230605791;#10;ip=64'd355030236726389;#10;ip=64'd529974940183956;#10;ip=64'd165370860002630;#10;ip=64'd337491883014368;#10;ip=64'd173955982213698;#10;ip=64'd212824546674804;#10;ip=64'd18357979033040;#10;ip=64'd396462137423370;#10;ip=64'd344489269643606;#10;ip=64'd331107488781342;#10;ip=64'd401332639464738;#10;ip=64'd32918101395946;#10;ip=64'd368104092918144;#10;ip=64'd160780840086408;#10;ip=64'd430089743062371;#10;ip=64'd157892017319667;#10;ip=64'd158462381610749;#10;ip=64'd123790118810293;#10;ip=64'd262879298977955;#10;ip=64'd529799286611159;#10;ip=64'd488233986223270;#10;ip=64'd547638321603475;#10;ip=64'd285131686687884;#10;ip=64'd556338120305653;#10;ip=64'd487143504771169;#10;ip=64'd431410597284617;#10;ip=64'd136253718959129;#10;ip=64'd400111089472257;#10;ip=64'd453476198141387;#10;ip=64'd276317542241782;#10;ip=64'd142237285888781;#10;ip=64'd113432275865793;#10;ip=64'd364520063516758;#10;ip=64'd125225213460866;#10;ip=64'd124344707468401;#10;ip=64'd294396567401905;#10;ip=64'd176790737993716;#10;ip=64'd216808838630653;#10;ip=64'd397750151505066;#10;ip=64'd26373057130794;#10;ip=64'd496488686770919;#10;ip=64'd267587062770538;#10;ip=64'd131737955785443;#10;ip=64'd558990543321844;#10;ip=64'd77619145636591;#10;ip=64'd559042476645382;#10;ip=64'd386430493134436;#10;ip=64'd448959511799118;#10;ip=64'd359033414943831;#10;ip=64'd409732629430972;#10;ip=64'd141381804210582;#10;ip=64'd393701708664165;#10;ip=64'd42263728504789;#10;ip=64'd395530023832103;#10;ip=64'd46185356083639;#10;ip=64'd293362744492551;#10;ip=64'd331460939645081;#10;ip=64'd355136654355101;#10;ip=64'd416986881512635;#10;ip=64'd296612941718408;#10;ip=64'd488997478224862;#10;ip=64'd226578471643146;#10;ip=64'd73314892719540;#10;ip=64'd237923758070672;#10;ip=64'd216608720732157;#10;ip=64'd520659018642157;#10;ip=64'd105437751572126;#10;ip=64'd188350034521574;#10;ip=64'd136207779748956;#10;ip=64'd13120397694442;#10;ip=64'd353195335000211;#10;ip=64'd238315824176265;#10;ip=64'd363609439811671;#10;ip=64'd520413272606668;#10;ip=64'd158844359173467;#10;ip=64'd88928460761659;#10;ip=64'd397283937120296;#10;ip=64'd560612815374967;#10;ip=64'd239279457113591;#10;ip=64'd386861906585659;#10;ip=64'd271741549290019;#10;ip=64'd343806775222642;#10;ip=64'd480645826376413;#10;ip=64'd327790109512732;#10;ip=64'd33603021914168;#10;ip=64'd527112388037717;#10;ip=64'd214484265098261;#10;ip=64'd411052416370110;#10;
        ip=64'd501838090752862;#10;ip=64'd330330296705262;#10;ip=64'd118557384101569;#10;ip=64'd208900462486969;#10;ip=64'd165298364833943;#10;ip=64'd536224056335022;#10;ip=64'd447732866271785;#10;ip=64'd184389579772140;#10;ip=64'd233608854663514;#10;ip=64'd81069391219868;#10;ip=64'd294864920049245;#10;ip=64'd163735403752189;#10;ip=64'd341197488271169;#10;ip=64'd1820706162357;#10;ip=64'd546631816644937;#10;ip=64'd370838913490358;#10;ip=64'd109032065371375;#10;ip=64'd339964427862925;#10;ip=64'd106721832160894;#10;ip=64'd334708161549928;#10;ip=64'd275894785247503;#10;ip=64'd77833700866251;#10;ip=64'd267501591283218;#10;ip=64'd295099737954661;#10;ip=64'd95432098993538;#10;ip=64'd507409126816274;#10;ip=64'd538333189599311;#10;ip=64'd224944992118647;#10;ip=64'd42370433743345;#10;ip=64'd509268740591107;#10;ip=64'd14683605271982;#10;ip=64'd468474941260401;#10;ip=64'd38347485134368;#10;ip=64'd26561871989463;#10;ip=64'd552184092749252;#10;ip=64'd511366878950980;#10;ip=64'd42431573537155;#10;ip=64'd307344291561581;#10;ip=64'd1576556301755;#10;ip=64'd120106765456840;#10;ip=64'd276722857333502;#10;ip=64'd397035470070311;#10;ip=64'd88009017645011;#10;ip=64'd471280708205467;#10;ip=64'd538118150510448;#10;ip=64'd496373666898978;#10;ip=64'd251330126428705;#10;ip=64'd31493391550982;#10;ip=64'd418492779197488;#10;ip=64'd168435287143829;#10;ip=64'd320869426607268;#10;ip=64'd19822938387106;#10;ip=64'd258816229632222;#10;ip=64'd359617340897220;#10;ip=64'd158501851288543;#10;ip=64'd295781677877933;#10;ip=64'd100512907323628;#10;ip=64'd355223285232519;#10;ip=64'd431410940073034;#10;ip=64'd500359767529111;#10;ip=64'd314774126365632;#10;ip=64'd474615360402726;#10;ip=64'd422043519146019;#10;ip=64'd19324793159674;#10;ip=64'd288560068613616;#10;ip=64'd102931122494764;#10;ip=64'd49714834719737;#10;ip=64'd353538945880083;#10;ip=64'd279645029040879;#10;ip=64'd536208458688175;#10;ip=64'd76371056564253;#10;ip=64'd268962943248816;#10;ip=64'd164198260155259;#10;ip=64'd475859662850135;#10;ip=64'd558309923703000;#10;ip=64'd13759158246199;#10;ip=64'd104352622724634;#10;ip=64'd383117154307607;#10;ip=64'd50981932789996;#10;ip=64'd531870023760703;#10;ip=64'd447085898932860;#10;ip=64'd560136302379470;#10;ip=64'd173753736557567;#10;ip=64'd328600618360733;#10;ip=64'd45840637514493;#10;ip=64'd248848268576596;#10;ip=64'd148256459775437;#10;ip=64'd541389968914834;#10;ip=64'd315250822385070;#10;ip=64'd268562700657170;#10;ip=64'd557831124666086;#10;ip=64'd236672333422075;#10;ip=64'd283252929074071;#10;ip=64'd518712588039529;#10;ip=64'd165875209940166;#10;ip=64'd425160092072958;#10;ip=64'd529441125772723;#10;ip=64'd89092489407613;#10;ip=64'd104018847974405;#10;ip=64'd265982174645724;#10;
        ip=64'd22900905150618;#10;ip=64'd279013968553980;#10;ip=64'd506778485091601;#10;ip=64'd498074249493987;#10;ip=64'd525275090717985;#10;ip=64'd2395564277545;#10;ip=64'd383626344055422;#10;ip=64'd194921149266529;#10;ip=64'd53492800965668;#10;ip=64'd386950813080721;#10;ip=64'd66299527442260;#10;ip=64'd386114941885516;#10;ip=64'd456080232519934;#10;ip=64'd495672003047972;#10;ip=64'd222943331040629;#10;ip=64'd237451177703722;#10;ip=64'd276340441460715;#10;ip=64'd449474748593781;#10;ip=64'd37581415565221;#10;ip=64'd539482192035200;#10;ip=64'd297250484140562;#10;ip=64'd197048493004545;#10;ip=64'd500818341914617;#10;ip=64'd188086129410107;#10;ip=64'd488008365966862;#10;ip=64'd149735573687976;#10;ip=64'd105622785933688;#10;ip=64'd143005856809599;#10;ip=64'd133578376039648;#10;ip=64'd76821898349613;#10;ip=64'd163920428965019;#10;ip=64'd227462424239368;#10;ip=64'd404271309778682;#10;ip=64'd488668432252242;#10;ip=64'd281619346458858;#10;ip=64'd298722796670245;#10;ip=64'd459125668492035;#10;ip=64'd315067066370578;#10;ip=64'd49724346763401;#10;ip=64'd445887743608892;#10;ip=64'd516198500720672;#10;ip=64'd38514289803191;#10;ip=64'd115417298589809;#10;ip=64'd532476041860658;#10;ip=64'd22444870178305;#10;ip=64'd171163571929812;#10;ip=64'd262995837633998;#10;ip=64'd188573913293368;#10;ip=64'd369081936445376;#10;ip=64'd544336935192010;#10;ip=64'd255862019330594;#10;ip=64'd559856665462458;#10;ip=64'd185140311517223;#10;ip=64'd398074817211298;#10;ip=64'd58008104825098;#10;ip=64'd307292053588251;#10;ip=64'd503002616323238;#10;ip=64'd101774565937304;#10;ip=64'd139366040569022;#10;ip=64'd398262289252141;#10;ip=64'd478958293458853;#10;ip=64'd176962861054670;#10;ip=64'd325633148986540;#10;ip=64'd164115801397488;#10;ip=64'd88654785009504;#10;ip=64'd63455893065089;#10;ip=64'd70795840110416;#10;ip=64'd556820404834619;#10;ip=64'd496252922463863;#10;ip=64'd187843877496782;#10;ip=64'd242443046864196;#10;ip=64'd51742573809393;#10;ip=64'd27103812516543;#10;ip=64'd128539952605923;#10;ip=64'd333969135484616;#10;ip=64'd541526362511105;#10;ip=64'd276981048416102;#10;ip=64'd537096545494302;#10;ip=64'd428504826116609;#10;ip=64'd34973926031242;#10;ip=64'd237344200705456;#10;ip=64'd233603747810312;#10;ip=64'd196477831630863;#10;ip=64'd158416574479184;#10;ip=64'd372004522954790;#10;ip=64'd437918593198043;#10;ip=64'd446372479279586;#10;ip=64'd294111542903923;#10;ip=64'd507749819918909;#10;ip=64'd482468793189330;#10;ip=64'd556689527676082;#10;ip=64'd450132335495005;#10;ip=64'd26561882652444;#10;ip=64'd511363003044467;#10;ip=64'd304481446309998;#10;ip=64'd66545818934060;#10;ip=64'd491921758108592;#10;ip=64'd40071431269444;#10;ip=64'd429521348543805;#10;ip=64'd109258372412341;#10;
        ip=64'd492117417398125;#10;ip=64'd116748245318213;#10;ip=64'd414546671529663;#10;ip=64'd95211636129804;#10;ip=64'd355777571607884;#10;ip=64'd198728568674203;#10;ip=64'd262403154671285;#10;ip=64'd424713725242829;#10;ip=64'd234705790721139;#10;ip=64'd56351196316496;#10;ip=64'd155546292451397;#10;ip=64'd477602932651908;#10;ip=64'd521176349274701;#10;ip=64'd433080764942472;#10;ip=64'd556639937396290;#10;ip=64'd410926970959868;#10;ip=64'd346209981831299;#10;ip=64'd288431278715030;#10;ip=64'd547134632315846;#10;ip=64'd328260011730876;#10;ip=64'd152101798498685;#10;ip=64'd163805088862870;#10;ip=64'd429744016648921;#10;ip=64'd123981466896196;#10;ip=64'd286242535699922;#10;ip=64'd98525385649523;#10;ip=64'd430051370556319;#10;ip=64'd399093414414436;#10;ip=64'd207332418328679;#10;ip=64'd141282175545293;#10;ip=64'd297915087977753;#10;ip=64'd220274033113130;#10;ip=64'd285661897457360;#10;ip=64'd478583804524434;#10;ip=64'd97067204352082;#10;ip=64'd255791766732058;#10;ip=64'd405927164550552;#10;ip=64'd61424768642389;#10;ip=64'd264684567887447;#10;ip=64'd327198612330874;#10;ip=64'd228026881833454;#10;ip=64'd105813686825780;#10;ip=64'd248502739474693;#10;ip=64'd441261855049594;#10;ip=64'd346223367408620;#10;ip=64'd53268602647886;#10;ip=64'd65124008148977;#10;ip=64'd486342245355864;#10;ip=64'd540739782616101;#10;ip=64'd58843520461460;#10;ip=64'd306391719098838;#10;ip=64'd15899941067785;#10;ip=64'd316060661804995;#10;ip=64'd495143730610215;#10;ip=64'd484158094684721;#10;ip=64'd488850162026480;#10;ip=64'd119317426746574;#10;ip=64'd284534174575553;#10;ip=64'd535025128249083;#10;ip=64'd372386161881462;#10;ip=64'd223262927435274;#10;ip=64'd236429879223797;#10;ip=64'd118873014498306;#10;ip=64'd9475800193741;#10;ip=64'd47425117938705;#10;ip=64'd524622827406086;#10;ip=64'd300424465406950;#10;ip=64'd229838788066287;#10;ip=64'd86862239278848;#10;ip=64'd184109066820780;#10;ip=64'd343787331887273;#10;ip=64'd518417084359855;#10;ip=64'd247731032002432;#10;ip=64'd494205601870100;#10;ip=64'd174214486983034;#10;ip=64'd186768788295859;#10;ip=64'd482207983314999;#10;ip=64'd158902192124152;#10;ip=64'd73457656383705;#10;ip=64'd18645183590998;#10;ip=64'd509894751192639;#10;ip=64'd153970337330873;#10;ip=64'd368653933246071;#10;ip=64'd213545348476355;#10;ip=64'd328219595331864;#10;ip=64'd174631310853266;#10;ip=64'd449174994711902;#10;ip=64'd506648197154482;#10;ip=64'd114255971201051;#10;ip=64'd77026160560810;#10;ip=64'd100985818747990;#10;ip=64'd364392881073848;#10;ip=64'd462091011955089;#10;ip=64'd437182973806886;#10;ip=64'd281401432690680;#10;ip=64'd315750284064961;#10;ip=64'd201832439835067;#10;ip=64'd483172845276324;#10;ip=64'd218158332323587;#10;ip=64'd385915276965347;#10;
        ip=64'd174552286324157;#10;ip=64'd197197859995996;#10;ip=64'd520261829177972;#10;ip=64'd154124630940652;#10;ip=64'd348345291947550;#10;ip=64'd268779044567477;#10;ip=64'd534359469218451;#10;ip=64'd316661087171691;#10;ip=64'd540970482935438;#10;ip=64'd283204753381961;#10;ip=64'd256202150667007;#10;ip=64'd377409600575216;#10;ip=64'd53140748496768;#10;ip=64'd62165338949555;#10;ip=64'd410186745194771;#10;ip=64'd58568372124543;#10;ip=64'd541423510656532;#10;ip=64'd160739964999512;#10;ip=64'd529651104706582;#10;ip=64'd59870610359031;#10;ip=64'd213447629726735;#10;ip=64'd342173193127989;#10;ip=64'd545190792560627;#10;ip=64'd303312973586569;#10;ip=64'd48723214881063;#10;ip=64'd263084961061495;#10;ip=64'd549888850563518;#10;ip=64'd35185953227819;#10;ip=64'd433852810391501;#10;ip=64'd24761890100966;#10;ip=64'd358882225027143;#10;ip=64'd547721783603707;#10;ip=64'd99954389985165;#10;ip=64'd2153660666090;#10;ip=64'd183870245785684;#10;ip=64'd184936924552048;#10;ip=64'd369881365422241;#10;ip=64'd388890177458544;#10;ip=64'd83430268637532;#10;ip=64'd202108860636669;#10;ip=64'd298170367232337;#10;ip=64'd64592670982912;#10;ip=64'd426289909384973;#10;ip=64'd289391640358689;#10;ip=64'd348662508320044;#10;ip=64'd506323485054029;#10;ip=64'd528684824095951;#10;ip=64'd276504679677249;#10;ip=64'd254080456609061;#10;ip=64'd126642047952945;#10;ip=64'd25377230139120;#10;ip=64'd438729773091090;#10;ip=64'd404006249676612;#10;ip=64'd178608993915853;#10;ip=64'd128251662002767;#10;ip=64'd436077237092060;#10;ip=64'd519656489051192;#10;ip=64'd394177913563735;#10;ip=64'd474632207876042;#10;ip=64'd261499928476941;#10;ip=64'd428418197368975;#10;ip=64'd127241376328602;#10;ip=64'd368350981243658;#10;ip=64'd342304374140833;#10;ip=64'd24122563409702;#10;ip=64'd270914300731571;#10;ip=64'd17646402661950;#10;ip=64'd479338312536756;#10;ip=64'd359428658750352;#10;ip=64'd217167284880929;#10;ip=64'd27459122596798;#10;ip=64'd5338696496932;#10;ip=64'd188424015829729;#10;ip=64'd53845604896642;#10;ip=64'd59487439194532;#10;ip=64'd227557051141650;#10;ip=64'd258997520644905;#10;ip=64'd534008991599462;#10;ip=64'd305381245486008;#10;ip=64'd490442432086665;#10;ip=64'd159150237849117;#10;ip=64'd533709242559454;#10;ip=64'd98925305078066;#10;ip=64'd239379486244956;#10;ip=64'd38264924496610;#10;ip=64'd398764326288835;#10;ip=64'd96817194993075;#10;ip=64'd518432687769212;#10;ip=64'd274255297854113;#10;ip=64'd486544622271597;#10;ip=64'd133845591971035;#10;ip=64'd466370211536413;#10;ip=64'd487434400044131;#10;ip=64'd175372619286803;#10;ip=64'd401132934169509;#10;ip=64'd45553957577854;#10;ip=64'd460313457139138;#10;ip=64'd115882983656728;#10;ip=64'd417759344338596;#10;ip=64'd85555240663755;#10;
        ip=64'd134209288230798;#10;ip=64'd236252579557749;#10;ip=64'd50654635426848;#10;ip=64'd387078452950102;#10;ip=64'd496619116565659;#10;ip=64'd450781451830972;#10;ip=64'd24683372396676;#10;ip=64'd403022236998396;#10;ip=64'd463536303335402;#10;ip=64'd287404561773493;#10;ip=64'd338241159784602;#10;ip=64'd546561332580057;#10;ip=64'd411468362064196;#10;ip=64'd473226910821451;#10;ip=64'd419793570846491;#10;ip=64'd430281078539833;#10;ip=64'd445275803377469;#10;ip=64'd234677632061946;#10;ip=64'd329434123739828;#10;ip=64'd514394512805837;#10;ip=64'd164050206491349;#10;ip=64'd353865931785966;#10;ip=64'd156624035938144;#10;ip=64'd211568532568807;#10;ip=64'd475006035187241;#10;ip=64'd498007335015799;#10;ip=64'd77733086056114;#10;ip=64'd535644164295210;#10;ip=64'd38728927281164;#10;ip=64'd460211644105777;#10;ip=64'd493382901194092;#10;ip=64'd48259660580174;#10;ip=64'd250749309205382;#10;ip=64'd34376208986091;#10;ip=64'd396963632978072;#10;ip=64'd333064034135419;#10;ip=64'd105600402298823;#10;ip=64'd91477433484584;#10;ip=64'd203850671211563;#10;ip=64'd168784874718009;#10;ip=64'd174331206638181;#10;ip=64'd514360685344896;#10;ip=64'd81213296146101;#10;ip=64'd511415691784083;#10;ip=64'd373010965981321;#10;ip=64'd97173641745402;#10;ip=64'd12927620480281;#10;ip=64'd270476772076226;#10;ip=64'd487623645653217;#10;ip=64'd205123366428936;#10;ip=64'd77004911781557;#10;ip=64'd115116717688229;#10;ip=64'd316728684858246;#10;ip=64'd550648197027569;#10;ip=64'd14273796260672;#10;ip=64'd433328329815736;#10;ip=64'd117341896382257;#10;ip=64'd114665609469341;#10;ip=64'd436091705783041;#10;ip=64'd111362462555076;#10;ip=64'd507548243812652;#10;ip=64'd341556118071111;#10;ip=64'd117982299070662;#10;ip=64'd341367296778284;#10;ip=64'd79284133915415;#10;ip=64'd489839563578476;#10;ip=64'd343316716562111;#10;ip=64'd510351447079436;#10;ip=64'd123053339909491;#10;ip=64'd15906690040338;#10;ip=64'd63708532109676;#10;ip=64'd374395174653859;#10;ip=64'd165656758489780;#10;ip=64'd115061474212145;#10;ip=64'd359567265588665;#10;ip=64'd231895682000110;#10;ip=64'd406102481131709;#10;ip=64'd436340644995578;#10;ip=64'd528451277816475;#10;ip=64'd82324803369168;#10;ip=64'd7406785540623;#10;ip=64'd186260256059584;#10;ip=64'd87956378439790;#10;ip=64'd509479945430089;#10;ip=64'd261022775022749;#10;ip=64'd548237177441683;#10;ip=64'd15430924760239;#10;ip=64'd355554883543477;#10;ip=64'd357362366589442;#10;ip=64'd15082504369846;#10;ip=64'd387682357482680;#10;ip=64'd124301027183705;#10;ip=64'd338775006812558;#10;ip=64'd502201227749636;#10;ip=64'd243480463189749;#10;ip=64'd228193433758368;#10;ip=64'd179532839909781;#10;ip=64'd14379955686134;#10;ip=64'd81910853594164;#10;ip=64'd465751075901815;#10;
        ip=64'd348713393416971;#10;ip=64'd236997304905458;#10;ip=64'd39589546421648;#10;ip=64'd497031556589966;#10;ip=64'd394303523291746;#10;ip=64'd457825575225945;#10;ip=64'd329214610077956;#10;ip=64'd532472393255943;#10;ip=64'd11991602296698;#10;ip=64'd83230235324806;#10;ip=64'd533531670172092;#10;ip=64'd404172096086643;#10;ip=64'd522306028688772;#10;ip=64'd27671413040236;#10;ip=64'd283701366772195;#10;ip=64'd440447729078619;#10;ip=64'd545856393818636;#10;ip=64'd57481137042691;#10;ip=64'd75082372920265;#10;ip=64'd249362419433125;#10;ip=64'd542501684481602;#10;ip=64'd68896596124547;#10;ip=64'd535749887111126;#10;ip=64'd163503989804318;#10;ip=64'd231705839194594;#10;ip=64'd485493211062017;#10;ip=64'd524774436413764;#10;ip=64'd215846335543972;#10;ip=64'd63276369767085;#10;ip=64'd295842610908245;#10;ip=64'd414261903459034;#10;ip=64'd266484911338005;#10;ip=64'd95520629296704;#10;ip=64'd451118345987462;#10;ip=64'd329309147068195;#10;ip=64'd245369563248269;#10;ip=64'd394393356736620;#10;ip=64'd120133254423146;#10;ip=64'd517963543652748;#10;ip=64'd383468866258786;#10;ip=64'd419052426090249;#10;ip=64'd198671439392472;#10;ip=64'd349522598702669;#10;ip=64'd509602147115657;#10;ip=64'd362069270271627;#10;ip=64'd443781264158562;#10;ip=64'd22303118797095;#10;ip=64'd260428022705942;#10;ip=64'd15853461610300;#10;ip=64'd479393589213688;#10;ip=64'd419778902580244;#10;ip=64'd337704128358101;#10;ip=64'd367402851108816;#10;ip=64'd83530409240506;#10;ip=64'd97061427163252;#10;ip=64'd219386734362160;#10;ip=64'd300214363147725;#10;ip=64'd240764593680882;#10;ip=64'd476888388291459;#10;ip=64'd466365365312505;#10;ip=64'd327488562606831;#10;ip=64'd520809344810386;#10;ip=64'd73637518028811;#10;ip=64'd179398335231127;#10;ip=64'd336511090000182;#10;ip=64'd224774825328810;#10;ip=64'd35013705236650;#10;ip=64'd237981848824794;#10;ip=64'd313720310144428;#10;ip=64'd402801478218905;#10;ip=64'd174896560893610;#10;ip=64'd92521474258207;#10;ip=64'd178433177773317;#10;ip=64'd35835484520801;#10;ip=64'd527621263708028;#10;ip=64'd286372497115081;#10;ip=64'd195025379170055;#10;ip=64'd379539077808192;#10;ip=64'd449901317243160;#10;ip=64'd35836911957793;#10;ip=64'd360405526771777;#10;ip=64'd175965627104994;#10;ip=64'd365342701128155;#10;ip=64'd201703696190484;#10;ip=64'd43699855218273;#10;ip=64'd157957598084265;#10;ip=64'd428533277124792;#10;ip=64'd30775472901661;#10;ip=64'd57004154492132;#10;ip=64'd338413139373411;#10;ip=64'd215567306895364;#10;ip=64'd193467404322766;#10;ip=64'd205657956351599;#10;ip=64'd74854694570884;#10;ip=64'd411538109269767;#10;ip=64'd258974282032069;#10;ip=64'd80056317298282;#10;ip=64'd369312257034699;#10;ip=64'd36042081121618;#10;ip=64'd48628156115854;#10;
        ip=64'd384623600661442;#10;ip=64'd406957034942134;#10;ip=64'd140725145290688;#10;ip=64'd154269622270305;#10;ip=64'd411914417216084;#10;ip=64'd435539108727611;#10;ip=64'd412278474797506;#10;ip=64'd345401394396629;#10;ip=64'd548087190342267;#10;ip=64'd558098316308587;#10;ip=64'd315481508535969;#10;ip=64'd106222639447539;#10;ip=64'd310770554102034;#10;ip=64'd417974884386986;#10;ip=64'd527494795130929;#10;ip=64'd281155256671197;#10;ip=64'd68774467816677;#10;ip=64'd432905456356026;#10;ip=64'd142780627919088;#10;ip=64'd550920554353665;#10;ip=64'd176332594611581;#10;ip=64'd253693085725395;#10;ip=64'd466003860181785;#10;ip=64'd196077520797913;#10;ip=64'd15786991190701;#10;ip=64'd474591960329046;#10;ip=64'd392573900139836;#10;ip=64'd358620206810363;#10;ip=64'd128610250685442;#10;ip=64'd147918700523519;#10;ip=64'd54894826961621;#10;ip=64'd185079718368601;#10;ip=64'd221877447282267;#10;ip=64'd464941392852971;#10;ip=64'd546970233553651;#10;ip=64'd425816575818336;#10;ip=64'd175299501782216;#10;ip=64'd112196519771999;#10;ip=64'd424625032429422;#10;ip=64'd371504019819394;#10;ip=64'd490630364192486;#10;ip=64'd202958854194653;#10;ip=64'd467417751397296;#10;ip=64'd398113819533258;#10;ip=64'd107318383125401;#10;ip=64'd360235590551131;#10;ip=64'd555207386200847;#10;ip=64'd396609442051770;#10;ip=64'd383613222621339;#10;ip=64'd376063174476632;#10;ip=64'd87483353397099;#10;ip=64'd270799347032251;#10;ip=64'd309130946476892;#10;ip=64'd88815363154102;#10;ip=64'd88162519262496;#10;ip=64'd475521547232526;#10;ip=64'd201197316152051;#10;ip=64'd293813977965301;#10;ip=64'd287317097932842;#10;ip=64'd9928624994278;#10;ip=64'd550344496254704;#10;ip=64'd99475141304812;#10;ip=64'd258032812671457;#10;ip=64'd328505985667717;#10;ip=64'd277560128615236;#10;ip=64'd486214125089126;#10;ip=64'd298386337215768;#10;ip=64'd77515919299748;#10;ip=64'd185332802632606;#10;ip=64'd358826373404061;#10;ip=64'd182698396088896;#10;ip=64'd55854138364545;#10;ip=64'd4395631879168;#10;ip=64'd43767118746026;#10;ip=64'd437085894433918;#10;ip=64'd509096205467757;#10;ip=64'd24282695177375;#10;ip=64'd489018023178684;#10;ip=64'd105784467650475;#10;ip=64'd361116089519808;#10;ip=64'd189149094217994;#10;ip=64'd547962074210876;#10;ip=64'd357863091409569;#10;ip=64'd307631027494673;#10;ip=64'd173716720652076;#10;ip=64'd517292292782125;#10;ip=64'd212444615948861;#10;ip=64'd213941868718524;#10;ip=64'd536613882349819;#10;ip=64'd345411902150087;#10;ip=64'd153092165511634;#10;ip=64'd75430665732431;#10;ip=64'd499066130260853;#10;ip=64'd166972840877860;#10;ip=64'd468185702217851;#10;ip=64'd479246038275046;#10;ip=64'd145445569891880;#10;ip=64'd358738312103304;#10;ip=64'd505254272953678;#10;
        $finish;
    end

endmodule
